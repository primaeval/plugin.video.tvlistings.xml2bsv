BBC1|1463874900|Weather for the Week Ahead|||0|0|Weather|
BBC1|1463875200|BBC News|21/05/2016||0|0|News|
BBC1|1463893200|Breakfast|||0|0|General Social,Political Issues,Economics|A round-up of national and international news, plus sports reports, weather forecasts and arts and entertainment features.
BBC1|1463901900|Match of the Day|Match of the Day - 2016 FA Cup Final Highlights||0|0|Football,Soccer|Crystal Palace v Manchester United. Action from the showpiece occasion at Wembley Stadium, along with post-match interviews and analysis. This was a repeat of the 1990 final, with current Palace boss Alan Pardew aiming to atone for being a member of the side that lost to United in a replay after the initial tie ended 3-3.
BBC1|1463904000|The Andrew Marr Show|22/05/2016||0|0|General News,Current Affairs|The political journalist presents a round-up of the week's stories, interviewing key figures and leafing through the Sunday papers.
BBC1|1463907600|The Big Questions|||9|17|Discussion,Debate|Nicky Campbell presents moral and religious discussions on topical issues from Wychwood School, Oxford.
BBC1|1463911200|Sunday Politics|22/05/2016||0|0|News Magazine,Current Affairs|The week's events at Westminster, presented by Andrew Neil. Including news and a regional round-up.
BBC1|1463915700|Bargain Hunt|Hay-on-Wye 19||40|16|Antiques,Collectibles|Tim Wonnacott presents the competition from Hay-on-Wye, Powys, where teams are guided by experts Charles Hanson and Jonathan Pratt through plenty of highs and lows. Meanwhile, the presenter stumbles across an interesting find with a well-travelled past.
BBC1|1463918400|BBC News|22/05/2016||0|0|National News|
BBC1|1463919000|Weather for the Week Ahead|||0|0|Weather|
BBC1|1463919300|Homes Under the Hammer|||0|0|Property|Martin Roberts and Lucy Alexander visit a flat in Stratford, east London and a semi-detached property in Whickham near Gateshead. The pair follow each lot to auction, and meet the people who bought them, before returning later to review the new owners' progress.
BBC1|1463921100|Escape to the Country|Herefordshire||12|40|Property|Nicki Chapman helps two Naval officers find their dream home in Herefordshire, but they cannot decide whether to increase their budget to more than £450,000. The presenter also joins in with the marigold harvest at a local organic farm.
BBC1|1463923800|Lose Weight for Love|Phil & Becky||1|1|Medicine,Health|Clinical psychologist Professor Tanya Byron and her team help couples who are locked in a cycle of over-eating, and are consequently threatening both their health and their relationship. In the first edition, cameras follow Becky and her partner Phil as they are separated for ten weeks in a bid to change their habits.
BBC1|1463927400|Nature's Epic Journeys|Caribou||1|2|Nature,Animals|Documentary following 100,000 caribou as they face bears, wolves, frozen rivers and rugged mountains to undertake the world's longest land migration. Liz Bonnin and a team of scientists track the herd as they travel 5,000km through the Arctic wilderness of Canada and Alaska, revealing insights into the lives of individual animals as they attempt the epic journey. Cameras capture the caribou as they fight to reach their calving grounds before they give birth - failure would spell disaster.
BBC1|1463931000|Lifeline|Church Housing Trust||0|0|General Education,Science|Julia Bradbury presents an appeal on behalf of Church Housing Trust, a charity that provides support for homeless people, and meets volunteers who were once homeless themselves.
BBC1|1463931600|Points of View|||0|0|General Education,Science|Jeremy Vine presents viewers' opinions on BBC shows and behind-the-scenes reports on new programmes.
BBC1|1463932500|Songs of Praise|||0|0|Folk,Traditional Music|A special episode for Dementia Awareness Week, in which Pam Rhodes discovers how a 1950s street has been recreated to help people with the condition. Plus, a pageant in Liverpool.
BBC1|1463934600|RHS Chelsea Flower Show 2016|||1|1|Gardening|New series. Sophie Raworth and Joe Swift present the first episode of this year's coverage from the Royal Horticultural Society's prestigious annual showcase, providing a look behind the scenes on the day before the showground officially opens to the public. Sophie and Joe discover how it takes three weeks of hard work to get everything ready for this week's grand opening, as well as providing a sneak preview of some of the spectacular gardens and exhibits set to make a big impression when the show gets underway.
BBC1|1463938200|BBC News|22/05/2016||0|0|National News|
BBC1|1463939400|BBC Regional News; Weather|22/05/2016||0|0|Regional News|
BBC1|1463940000|Countryfile|Veggie Theme||0|0|Nature,Animals|A special episode for National Vegetarian Week, in which Matt Baker visits Jersey during the royal potato harvest and Ellie Harrison creates a landscape photograph with vegetables. Naomi Wilkinson samples some Indian vegetarian recipes, sheep farmer Gareth Wyn Jones and free runner Tim Shieff debate the pros and cons of veganism, and Adam Henson visits an underground urban farm. Plus, Tom Heap investigates why many vegetable growers face going out of business. Including Weather For The Week Ahead.
BBC1|1463943600|Antiques Roadshow|Tredegar House 1||37|9|Antiques,Collectibles|Fiona Bruce and the team visit Tredegar House near Newport in Wales, where members of the public bring along treasured antiques and collectibles. Items of interest include a tapestry woven in tribute to Status Quo, a carved coconut steeped in 18th-century maritime history and a frog-shaped brooch. A former Mastermind champion shows off the glass vase he won, and a Second World War veteran tells the story of a daring mission to inspect German defences before the D-Day landings - and how he came to have a packet of cigarettes from Field Marshal Rommel.
BBC1|1463947200|Wallander|The White Lioness||4|1|General Movie,Drama|New series. Kenneth Branagh stars as the world-weary Swedish detective in a fourth and final series of adaptations of Henning Mankell's novels. Wallander travels to Cape Town to investigate the disappearance of a Swedish woman. He uncovers a complex conspiracy behind the mystery, and is also confronted with a nation that has reached a turning point in its history.
BBC1|1463952600|BBC News|22/05/2016||0|0|National News|
BBC1|1463953800|BBC Regional News; Weather|22/05/2016||0|0|Regional News|
BBC1|1463954400|Room 101 - Extra Storage|||4|5|Comedy|An extended edition of the show in which chat-show host Jonathan Ross, former England cricket captain Michael Vaughan and comedienne Sara Pascoe tell Frank Skinner what really gets on their wick. The celebrities' gripes include pick 'n' mix, misuse of the word `literally' and the Grim Reaper.
BBC1|1463956800|Athletics|Athletics: Diamond League Rabat Highlights||0|0|Athletics|Gabby Logan presents action from the third Diamond League event of the season, held at Prince Moulay Abdellah Stadium in Rabat, Morocco.
BBC1|1463960400|Weather for the Week Ahead|||0|0|Weather|
BBC1|1463960700|BBC News|22/05/2016||0|0|News|
BBC1|1463979600|Breakfast|||0|0|General Social,Political Issues,Economics|Round-up of national and international news, plus the latest from the money markets.
BBC1|1463991300|Council House Crackdown|||2|1|General Education,Science|New series. The return of the programme that follows local authority housing officers as they track down social housing cheats, beginning with Croydon Council investigating a fraudulent tenant. Luke Doonan and Michelle Ackerley present.
BBC1|1463994000|Homes Under the Hammer|||19|50|Property|Lucy Alexander, Martin Roberts and Dion Dublin meet investors who have bought properties in Doncaster, the Kent town of Strood and High Hatton in Shropshire.
BBC1|1463997600|Family Finders|||0|0|General Education,Science|New series. The work of Britain's ever-growing army of commercial tracing companies and independent genealogy detective agencies. Together with more established bodies such as the Salvation Army, these dedicated staff devote their time to tracking down and reuniting lost family members.
BBC1|1464000300|Break-in Britain - The Crackdown|Getaway Bus||2|1|General Education,Science|Police investigate a burglary at the Leeds home of pensioners Nick and Avril, where Keeley sets out to improve the couple's security, and Dan goes to the aid of a South Wales woman whose house has been ransacked.
BBC1|1464002100|Bargain Hunt|Westpoint 17||44|0|Antiques,Collectibles|Paul Laidlaw presents from the Westpoint Arena in Exeter as experts Richard Madley and Charlie Ross help two teams to make the most profit at auction. Paul also visits the city's Met Office to learn about the history of weather forecasting.
BBC1|1464004800|BBC News at One; Weather|23/05/2016||0|0|News|
BBC1|1464006600|BBC Regional News and Weather|||0|0|Regional News|
BBC1|1464007500|Doctors|The Collector||18|35|Soap,Melodrama|Jimmi visits Mrs Tembe and uncovers her issues, while Karen is stressed by a home visit by her social worker and Emma has to deal with a policeman accused of theft.
BBC1|1464009300|For What It's Worth|||2|1|Antiques,Collectibles|New series. Fern Britton returns with the game show in which three pairs of contestants try to amass a valuable collection of antiques and collectibles by answering general knowledge questions, with the value of the items they win being converted to a cash prize. With expert advice from Charlie Ross.
BBC1|1464012000|Escape to the Country|Oxfordshire||16|61|Property|Jules Hudson is on a property hunting mission in Oxfordshire with two newlyweds who have £400,000 to spend in an attempt to return to their rural roots and start a family. Jules also visits a bespoke bookbinder keeping traditional, handcrafted techniques alive.
BBC1|1464014700|RHS Chelsea Flower Show 2016|||1|2|Gardening|Nicki Chapman and James Wong take the first official look at the Royal Horticultural Society's show, which opened its gates to the world at 6.30am, with Carol Klein in the Great Pavilion to take a closer look at life-changing plants and ex-footballer Sol Campbell shares his love of gardening. The team captures all the buzz as celebrities and VIPs take their first look and reports on how Chelsea is preparing for the arrival of the Queen.
BBC1|1464017400|Flog It|Dorset 21||13|29|Antiques,Collectibles|Antiques experts Catherine Southon and Mark Stacey value items and collectibles brought in by the public to Lulworth Castle in Dorset. Plus, presenter Paul Martin explores the turbulent history of the Weld family and the anti-Catholic persecution they were subject to for more than 300 years.
BBC1|1464020100|Pointless|||15|24|Quiz Show|Quiz show in which pairs of contestants try to score the fewest points possible by giving the least obvious correct answers to questions posed to 100 people before the show. At the end of each round, the team with the most points is eliminated until the final two pairs battle for the chance to compete for a cash prize. Presented by Alexander Armstrong and Richard Osman.
BBC1|1464022800|BBC News at Six; Weather|23/05/2016||0|0|News|
BBC1|1464024600|BBC Regional News Programmes|||0|0|Regional News|
BBC1|1464026100|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Vote Leave campaign.
BBC1|1464026400|The One Show|23/05/2016||0|0|General Education,Science|The first visit of the week to the One Show studio, where Matt Baker and Alex Jones present the usual mix of topical stories and celebrity chat.
BBC1|1464028200|RHS Chelsea Flower Show 2016|||1|3|Gardening|Sophie Raworth and Joe Swift present coverage of the horticultural event from around the showground, including footage from the Queen's annual visit. Meanwhile, the Chelsea team guides viewers through show-stopping gardens and exhibits.
BBC1|1464030000|EastEnders|||0|0|Soap,Melodrama|All hell breaks loose for the Beales when Bobby strikes again, leaving Jane fighting for her life - and as if that weren't bad enough, the troubled youngster then announces what he has just done to the assembled guests at Stacey and Martin's wedding party. Can Ian continue to protect his son under such shocking circumstances? Meanwhile, Roxy comes looking for Amy at the Vic, where Linda tries to get her to open up about Dean, and Jack Ronnie spots Andy fleeing the Square.
BBC1|1464031800|Panorama|Antibiotic Crisis - Panorama||0|0|Documentary|Tom Heap reports on how resistance to prescribed antibiotics could become a serious public health threat. He also investigates how antibiotics used in farming could lead to a rise in superbugs and meets patients who have found the drugs they have been prescribed have no effect.
BBC1|1464033600|Peter Kay's Comedy Shuffle|||1|6|Comedy|A final selection from the career of the comedian, actor, writer and director, featuring Peter appearing with Catherine Tate's Nan as well as his observations on family weddings and more of Max and Paddy's misadventures. Last in the series.
BBC1|1464035400|I Want My Wife Back|||1|6|Sitcom|Murray drops one of Bex's dresses round to her at Keeley's flat for her parents' anniversary party that evening and finds a positive pregnancy test in her temporary bedroom, prompting him to try everything he can do to get her back. At the bank, he tries to get a definitive answer from Emma on whether or not anything happened between them that night, but she is distracted and unable to give him a straight answer, while Keeley has a big decision about the future of her relationship. Comedy, starring Ben Miller and Caroline Catz. Last in the series.
BBC1|1464037200|BBC News at Ten|23/05/2016||0|0|News|
BBC1|1464039000|BBC Regional News and Weather|||0|0|Regional News|
BBC1|1464039900|Have I Got a Bit More News for You|||51|7|Comedy|Gary Lineker hosts an extended edition of the satirical quiz, with panellists Ross Noble and Samira Ahmed joining team captains Ian Hislop and Paul Merton.
BBC1|1464042600|The Graham Norton Show|||19|9|Comedy|Hollywood stars Ryan Gosling and Russell Crowe talk about their new film The Nice Guys, while double Oscar-winner Jodie Foster promotes her directorial feature Money Monster. Plus, Elton John and Bright Light Bright Light, aka Rod Thomas, perform All in the Name. The host also subjects more audience members to the dreaded red chair - so their stories had better be good.
BBC1|1464045300|Weather for the Week Ahead|||0|0|Weather|
BBC1|1464045600|BBC News|23/05/2016||0|0|News|
BBC1|1464066000|Breakfast|||0|0|General Social,Political Issues,Economics|Round-up of national and international news, plus the latest from the money markets.(n)
BBC1|1464077700|Council House Crackdown|||2|2|General Education,Science|Michelle Ackerley follows the case of a grandmother who appears in court after illegally subletting her council flat, and an assignment involving a missing mother and daughter.(n)
BBC1|1464080400|Homes Under the Hammer|||19|51|Property|Lucy Alexander, Martin Roberts and Dion Dublin explore a semi in Chingford, London, a one-bedroom flat in Brighton and a Victorian terrace in Normanton, Derby.(n)
BBC1|1464084000|Family Finders|Belinda & Alex/Barb & Sybil||2|2|General Education,Science|Inspired by an old letter from a mysterious relative in Peru, Belinda O'Brien researches her family history, and Barbara Cohen attempts to finds out more about her own family.(n)
BBC1|1464086700|Break-in Britain - The Crackdown|Hunt for Gold||2|2|General Education,Science|Dan Donnelly makes a Leeds home secure, and police hope the burglar's dropped phone will help identify their man. Meanwhile, Keeley Donovan hunts for a Swansea motorbike thief.(n)
BBC1|1464088500|Bargain Hunt|Lincoln 1||41|1|Antiques,Collectibles|Mark Stacey and Natasha Raskin offer their expert opinions as two teams attempt to pick up bargains at the Lincolnshire Showground, where one friendship is pushed to the limit. Meanwhile, host Tim Wonnacott takes time out to visit one of the UK's finest Georgian houses.(n)
BBC1|1464091200|BBC News at One; Weather|24/05/2016||0|0|News|
BBC1|1464093000|BBC Regional News and Weather|||0|0|Regional News|
BBC1|1464093900|Doctors|Just Say No||18|36|Soap,Melodrama|Sid tries to persuade a university lecturer to stop taking drugs, Al reluctantly gives a presentation, and Heston is forced to consider the practical benefits of Ruhma's religion.(n)
BBC1|1464095700|For What It's Worth|||2|2|Antiques,Collectibles|Fern Britton hosts the game show in which three pairs of contestants try to amass a valuable collection of antiques and collectibles by answering general knowledge questions, with the value of the items they win being converted to a cash prize.(n)
BBC1|1464098400|Escape to the Country|North Yorkshire||13|47|Property|Alistair Appleton heads to North Yorkshire, where he helps a couple with a budget of £550,000 find a rural property suitable to let as a holiday home. The presenter also visits Whitby Folk Festival, an annual event that celebrates traditional music and dance from around the British Isles.(n)
BBC1|1464101100|RHS Chelsea Flower Show 2016|||1|5|Gardening|It's medals day at the annual event, so Nicki Chapman and James Wong join the judges early on to discover who has won what in the all-important handout. Bake Off supremo Mary Berry reveals that she knows her way around the garden as well the kitchen, and Kate Adie discusses her new-found passion for horticulture.(n)
BBC1|1464103800|Flog It|Margam Country Park||14|44|Antiques,Collectibles|Mark Stacey and Charles Hanson are in Margam Country Park in south Wales to value items brought in by the public, while presenter Paul Martin finds out about the link between the estate and the nearby Port Talbot steelworks.(n)
BBC1|1464106500|Pointless|||12|17|Quiz Show|Quiz show in which pairs of contestants try to score the fewest points possible by giving the least obvious correct answers to questions posed to 100 people before the show. At the end of each round, the team with the most points is eliminated until the final two pairs battle for the chance to compete for a cash prize. Presented by Alexander Armstrong and Richard Osman.(n)
BBC1|1464109200|BBC News at Six; Weather|24/05/2016||0|0|News|
BBC1|1464111000|BBC Regional News and Weather|||0|0|Regional News|
BBC1|1464112500|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|A referendum broadcast by the Stronger in Europe campaign, ahead of the Referendum on the United Kingdom's membership of the European Union, on June 23rd.(n)
BBC1|1464112800|The One Show|||0|0|General Education,Science|Another mix of nationwide reports and live studio-based chat, hosted by Matt Baker and Alex Jones.(n)
BBC1|1464114600|EastEnders|||0|0|Soap,Melodrama|Ian and his family wait anxiously at the hospital for news on Jane - except for Bobby, whose world is thrown into turmoil when he is arrested for the attack on his stepmother. Sharon tries to help her friends by taking control of the situation, although she is stunned by a turn of events, and a concerned Denise reaches out to an old friend.(n)
BBC1|1464116400|Holby City|When I Grow Up||18|33|General Movie,Drama|Arthur is determined to prove his worth in the face of Hanssen's ambitions, but he struggles to keep his personal and professional lives separate, leaving him forced to make a tough decision. Oliver sees a chance to get back together with Zosia, but ends up in need of Cara's support when he pushes things too far. Raf comes to see Naomi in a new light, and makes a personal sacrifice.(n)
BBC1|1464120000|In the Club|||2|4|General Movie,Drama|With Shelly keeping baby Sebastian with her on the ward overnight, an anxious Andrew and Nathan prepare to bring him home again. Andrew's convinced something's going to go wrong and that Shelly will change her mind, while Nathan struggles to keep him calm. But neither of them is prepared for the shock of what is waiting for them at the hospital. Meanwhile, Maxine's day is thrown into chaos when she gets a call from her husband Micky, saying he's on his way home, and things get increasingly complicated for Roanna as she and Ray continue to meet in secret.(n)
BBC1|1464123600|BBC News at Ten|24/05/2016||0|0|News|
BBC1|1464125400|BBC Regional News and Weather|||0|0|Regional News|
BBC1|1464126300|Last Whites of the East End|||0|0|General Education,Science|Newham in East London has the lowest white British population in the UK. This film tells the stories of the last caucasian Eastenders who have started to feel `like foreigners in their own land'. Through the journeys of people leaving, or staying in a place that no longer feels like home, cameras follow the last whites in Newham as the world changes around them.(n)
BBC1|1464129900|The Truth About|The Truth About Dementia||2|1|Medicine,Health|In the first of three documentaries focusing on health matters, Angela Rippon, who lost her mother to Alzheimer's, presents the latest scientific research about dementia - of which Alzheimer's is the most common form. She undergoes tests to see if she has any early signs, learns some surprising ways that may help prevent dementia and visits a number of people living with the disease. She also meets families that carry a gene for early onset Alzheimer's, discovering how they could be the best hope of finding a cure for this devastating disease.(n)
BBC2|1463874000|Elena||2011|0|0|General Movie,Drama|A woman from a poor background marries a richer man. However, when the husband becomes seriously ill, he announces his plan to cut her out of the will and bequeath everything to his daughter from a previous marriage, leaving her desperate to secure a stable future for herself and her son. Drama, starring Nadezhda Markina and Andrey Smirnov. In Russian.
BBC2|1463880000|This Is BBC Two|||0|0|General Show,Game Show|Preview of upcoming programmes from BBC Two.
BBC2|1463891700|The Great Chelsea Garden Challenge|The Final||1|4|Gardening|The three remaining competitors visit the RHS Headquarters in Wisley for the grand final of the garden design competition. Here, they are given five days - and their biggest budget yet - to put together showpiece gardens that will impress judges James Alexander-Sinclair and Ann-Marie Powell, and prove they are worthy of going to Chelsea. Joe Swift provides expert tips, with the winning designer earning the chance to put together a garden for the Main Avenue at RHS Chelsea Flower Show 2015. Last in the series.
BBC2|1463895300|This Farming Life|||1|10|General Education,Science|Sybil prepares for George's 50th birthday and the arrival of her sister and niece from England, while persistent rain means Martin's cattle are yet to be turned out of their winter sheds into the fields. Bobby and Anne hold an open day to educate the public about farming and John has to urgently call the vet when one of his heifers gets into difficulty calving.
BBC2|1463898900|Gardeners' World|||49|10|Gardening|Monty Don plants up containers to add colour to his jewel garden at Longmeadow. He also turns his attention to overcrowded ornamental grasses, which need to be split and replanted. Carol Klein takes a look at plants able to survive in cracks and crevices and gives her recommendations for garden plants that will thrive in similar conditions. Plus, Zephaniah Lindo takes a trip to Wales to meet a fellow primula enthusiast.
BBC2|1463900700|Countryfile|Countryfile Spring Special||0|0|Nature,Animals|The team reports on signs of spring around the country, with Ellie Harrison monitoring pods of returning dolphins in Cardigan Bay and John Craven visiting a hay meadow in Wiltshire that's uninterrupted agricultural history has created a rare environment that has lasted for more than 800 years. Matt meets a couple who have turned a Roman fort on Alderney into a bird observatory, while Anita Rani spends a day in with fishermen in Newlyn as they haul in lobster pots.
BBC2|1463904000|The Beechgrove Garden|||38|8|Gardening|Jim McColl tries out a range of gadgets for growing tomatoes as he starts off some new varieties, and he and George Anderson visit the world's largest cut-flower auction, at Aalsmeer near Amsterdam. Scone Palace head gardener Brian Cunningham continues his revamp of the alpine garden, finishing off the hard landscaping and starting the planting.
BBC2|1463905800|Saturday Kitchen Best Bites|||0|0|Cooking|James Martin presents highlights of the series, recalling his favourite moments from previous years in the kitchen. Featuring an archive programme presented by Rick Stein.
BBC2|1463911200|Live Athletics|Live Athletics: Great Manchester Run||0|0|Athletics|Jonathan Edwards presents coverage of the 14th staging of the event, as approximately 40,000 runners take part. Another stellar cast of athletes are set to be involved, including three-time Olympic gold medallist Tirunesh Dibaba, making her comeback in the women's elite race after time off to have a baby in 2015. With commentary by Steve Cram, Paula Radcliffe and Andrew Cotter, and reports from Denise Lewis and Phil Jones.
BBC2|1463918400|Custer of the West||1967|0|0|Biopic|Historical biopic based on the life of the American cavalry commander who achieved military success during the Civil War, and was sent to seize land for the US government, ultimately meeting his end at the Battle of the Little Bighorn. Starring Robert Shaw, Mary Ure, Jeffrey Hunter, Ty Hardin and Lawrence Tierney.
BBC2|1463926500|Flog It|Stockport 2||11|50|Antiques,Collectibles|Antiques experts Mark Stacey and Philip Serrell head to Stockport Town Hall in Greater Manchester to value the collectibles of members of the public, including a pair of charcoal drawings by artist Trevor Grimshaw and some gold European coins. Plus, presenter Paul Martin visits Manchester Art Gallery, where he admires the work of pre-Raphaelite painter Ford Madox Brown.
BBC2|1463929200|Swimming: European Championships|||0|0|Swimming|Helen Skelton presents live coverage of the final day of swimming events at the European Aquatics Championships, from the Aquatics Centre at Queen Elizabeth Olympic Park in London. Two years ago in Berlin, Team GB had a day to remember when Fran Halsall, Jazz Carlin and the men's 4x100m medley relay team all won gold in their respective events, with Great Britain topping the final medal table in the process.
BBC2|1463936400|Athletics|Athletics: Great Manchester Run Highlights||0|0|Athletics|Action from the 14th annual staging of the 10k race, as elite athletes and thousands of fun runners competed. With commentary by Steve Cram, Paula Radcliffe and Andrew Cotter.
BBC2|1463940000|Britain's Ultimate Pilots: Inside the RAF|||1|3|Documentary|The Red Arrows mark the end of an era as they appear in a succession of airshows, including events where they fly alongside a Vulcan bomber and a Chinook helicopter. The pilots have to undergo gruelling underwater training before they can appear at a planned display in Blackpool, but it seems that the performance may be grounded as a result of high winds.
BBC2|1463943600|World Cup 1966: Alfie's Boys|||0|0|Documentary|David Jason presents a documentary about how Alf Ramsey recruited the England football team that won the world cup in 1966, and was able to unite the members into a world class side. Featuring archive footage of the team in action and contributions from Bobby Charlton, Jack Charlton, Jimmy Greaves, George Cohen, Tina Moore, Harry Redknapp, Terry Venables, Geoff Hurst and Gordon Banks.
BBC2|1463949000|Horizon|Horizon: E-Cigarettes - Miracle or Menace?||0|0|Documentary|Michael Mosley investigates the dramatic rise in e-cigarettes in recent years, and questions whether they are a health risk or a better alternative to smoking. He reports on the content of e-cigarettes, meets scientists who are studying their effects and takes up vaping himself to see how it effects his health.
BBC2|1463952900|Stupid Man, Smart Phone|Norway||1|2|General Education,Science|Russell Kane travels through Norway, heading into the Arctic Circle in the hope of seeing the Northern Lights. He is accompanied on his journey by Youtube stars Rose and Rosie, and together they rely on a smartphone to provide answers to all the challenges the expedition throws their way.
BBC2|1463955900|Later - with Jools Holland|||48|5|General Music,Ballet,Dance|Extended edition of the music programme. Iggy Pop makes his debut on the show, performing tracks from his recent album Post Pop Depression, recorded with Josh Homme, who joins him on stage with fellow Queens of the Stone Age band member Dean Fertita and Arctic Monkeys drummer Matt Helders. Plus, performances by Lou Doillon, Protoje, Graham Nash, Blossoms and Margo Price.
BBC2|1463959800|Countryfile|Countryfile Spring Special||0|0|Nature,Animals|The team reports on signs of spring around the country, with Ellie Harrison monitoring pods of returning dolphins in Cardigan Bay and John Craven visiting a hay meadow in Wiltshire that's uninterrupted agricultural history has created a rare environment that has lasted for more than 800 years. Matt meets a couple who have turned a Roman fort on Alderney into a bird observatory, while Anita Rani spends a day in with fishermen in Newlyn as they haul in lobster pots.
BBC2|1463963100|Holby City|Running Out||18|32|General Movie,Drama|Zosia oversteps the mark and accuses a patient of a media leak, leaving Oliver with an unwelcome dilemma. As his suspicions spiral out of control, Zosia makes a gut-wrenching decision. Dominic faces his fears when he encounters someone with a painful past, and Serena returns to find Bernie helping out on AAU. However, her gratitude is short-lived when she discovers the real reason for the surgeon's presence on the ward.
BBC2|1463966700|This Is BBC Two|||0|0|General Show,Game Show|Preview of upcoming programmes from BBC Two.
BBC2|1463980500|Homes Under the Hammer|||20|12|Property|Dion Dublin, Martin Roberts and Lucy Alexander meet the new owners of an old barbershop in Rochdale, Lancashire, a bungalow in Alsager, Cheshire and a piece of land in Eccles, Kent. They reveal their ideas for redevelopment - but will everything go according to plan?.
BBC2|1463984100|Flog It|||0|0|Antiques,Collectibles|Paul Martin recalls trips to Muncaster Castle in Cumbria, the Bowes Museum in Co Durham, the Grand Pier in Weston-super-Mare in Somerset and Norwich Cathedral, where antiques experts inspected items ranging from an antique tipstaff to a piece of Bernard Leach pottery.
BBC2|1463986800|Food Detectives|||1|3|General Education,Science|Alice Roberts tests the claim that drinking artificially sweetened drinks encourage people to eat more than they would have done had they consumed a sugary drink, while Sean Fletcher investigates whether it is worth paying for a premium product when a money-saving basic alternative as just as good in terms of health and taste. Tom Kerridge heads in Glasgow to advise a viewer on preparing perfect Yorkshire puddings.
BBC2|1463988600|Gardeners' World|||49|9|Gardening|As the growing season gathers pace, Monty Don sows vegetables and plants out the scented plants he brought back from the Malvern Spring Festival. Carol Klein delves into the hedgerows and rooting at the bases of walls, fences and trees as she begins her journey to investigate why plants thrive in challenging conditions. The programme also returns to Sissinghurst, Kent, to learn about the changes head gardener Troy Scott-Smith is planning to Vita Sackville-West's 1930s creation.
BBC2|1463990400|Victoria Derbyshire|23/05/2016||0|0|News Magazine,Current Affairs|Daily news and current-affairs programme offering discussion of breaking stories, exclusive interviews and audience interaction via social media.
BBC2|1463997600|BBC Newsroom Live|23/05/2016||0|0|General News,Current Affairs|A chance to stay up to date on the day's leading stories, with the latest breaking news as it happens.
BBC2|1464001200|Daily Politics|23/05/2016||0|0|Discussion,Debate|Parliamentary proceedings interspersed with discussions, interviews and reports from correspondents around the country. Presented by Jo Coburn.
BBC2|1464004800|Athletics|Athletics: Diamond League Rabat Highlights||0|0|Athletics|Gabby Logan presents action from the third Diamond League event of the season, held at Prince Moulay Abdellah Stadium in Rabat, Morocco.
BBC2|1464008400|Paul Hollywood's Pies & Puds|||1|9|Cooking|The baker continues his exploration of British food by sampling a marshmallow company's products and their perfect accompaniments to his sticky toffee pudding. Plus, he shares his recipes for salted caramel coffee eclairs and picnic empanadas.
BBC2|1464010200|The TV That Made Me|Gok Wan||1|10|Popular Culture,Traditional Arts|Gok Wan joins Brian Conley to revisit some classic television series of his formative years. From the magic and mystery of Japanese children's drama Monkey, to the pan-European quiz show Going for Gold, via groundbreaking, anarchic pop series The Tube, these were the shows that apparently helped shape Gok into the style icon that he is today.
BBC2|1464012000|Holiday of My Lifetime with Len Goodman|Matt Allwright||1|11|Tourism,Travel|The Strictly Come Dancing judge takes consumer journalist Matt Allwright on a journey to Teignmouth and Shaldon in Devon, to recreate a family holiday experience from 1977. Among the activities on the pair's to-do list are mackerel fishing, arcade gaming on penny slot machines, and a trip to Babbacombe Model Village in nearby Torquay.
BBC2|1464014700|This World|The Tea Trail with Simon Reeve||0|0|General Education,Science|In the first of two This World documentaries examining the stories behind the nation's favourite beverages, adventurer and broadcaster Simon Reeve looks at the production of tea. He begins in the Kenyan coastal city of Mombasa, where most of the leaves for teabags are bought at auction, before travelling through eastern Africa to meet some of the millions of people who pick, pack and transport it. He drinks tea with everyone from Maasai cattle herders to the descendants of the original plantation owners, and hears claims of low wages and child labour.
BBC2|1464018300|Great British Railway Journeys|Manchester to Birkenhead||5|1|General Education,Science|Armed with a copy of George Bradshaw's Victorian Railway Guidebook, Michael Portillo embarks on another journey around the country to discover how the railways have affected people and communities, and the legacy they have left behind. He begins in Manchester, where he finds out how the world's first industrialised city produced a revolutionary political movement, and learns about the railway workers who founded one of the most successful football clubs of all time. Along the way, the presenter does the washing in Port Sunlight - a model village on the Wirral - and hears stories about the aptly named George Francis Train's time in Birkenhead, Merseyside.
BBC2|1464020100|Bargain Hunt|Deene Park 25||36|27|Antiques,Collectibles|Experts Kate Bateman and Thomas Plant head to Deene Park in Northamptonshire, where two teachers and a pair of murder mystery actors put their bargain-spotting abilities to the test. Meanwhile, Tim Wonnacott visits the Charterhouse School in Guildford, Surrey, which has produced some of Britain's finest musicians, including members of the pop group Genesis.
BBC2|1464022500|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Vote Leave campaign.
BBC2|1464022800|Eggheads|||17|59|Game Show,Quiz|Jeremy Vine hosts the quiz in which the winners of famous game shows including Mastermind and Who Wants to Be a Millionaire? work as a team to tackle a new set of challengers hoping to win a cash prize.
BBC2|1464024600|Countryfile Spring Diaries|New Life!||1|1|Rural,Agricultural|A look at the impact of the arrival of spring around the nation, with John Craven and Keeley Donovan kicking things off by investigating what makes the season's weather so special. Jules Hudson takes to the saddle to find out why this is a crucial time for New Forest ponies and Margherita Taylor reports on how to tap trees for silver birch sap. Every day this week, Paul Martin will be breathing new life into his Victorian smallholding in Wiltshire, starting with the hunt for a perfect breed of sheep to help restore his fields.
BBC2|1464026400|Antiques Road Trip|||0|0|Antiques,Collectibles|Christina Trevanion and Thomas Plant start their trip in north Wales, before travelling through Warwickshire and Essex in a 1962 Bedford van. On their way, they witness a spectacular Battle of Britain air show and head for the auction showdown in Winchcombe, Gloucestershire.
BBC2|1464030000|RHS Chelsea Flower Show 2016|||1|4|Gardening|Monty Don and Joe Swift present further coverage of the horticultural event, which has been held in the grounds of the Royal Hospital Chelsea since 1913. There are highlights of the Queen's annual visit and a look ahead to tomorrow's medals announcement as the presenters predict the designer they think will scoop the coveted best show garden award. Plus, actor Tom Hollander joins Monty and Joe to chat about his love of gardening.
BBC2|1464033600|The Great British Sewing Bee|||4|2|General Education,Science|Claudia Winkleman sets the remaining contestants three challenges designed to test different fabric handling skills on children's clothing.  Firstly, they must carefully follow a pattern to make baby grows from stretch cotton jersey and then show they can handle slippery satin and chiffon by transforming an adult bridesmaid's dress into a garment for a boy or a girl. Finally, they have to create perfectly fitted woollen capes, before judges Patrick Grant and Esme Young decide who leaves the competition.
BBC2|1464037200|Upstart Crow|The Apparel Proclaims the Man||1|3|Sitcom|Will hopes to move up in the world when he is invited to a high-society party hosted by Lord Southampton, but is unsure what a poorly-educated country boy should wear to one of London's most upmarket events. The playwright's rival Sir Robert Greene offers him some fashion tips, but is it a double bluff, a triple bluff, or something even more fiendish? Ben Elton's comedy about William Shakespeare's family and professional lives, starring David Mitchell as the Bard, with Mark Heap and Liza Tarbuck.
BBC2|1464039000|Newsnight|23/05/2016||0|0|News Magazine,Current Affairs|Analysis of the day's events, presented by Evan Davis.
BBC2|1464042600|Weather|||0|0|Weather|
BBC2|1464042900|Horizon|Curing Alzheimer's||0|0|Documentary|Documentary investigating scientific breakthroughs in research on Alzheimer's disease, which are bringing hope to millions of sufferers across the world. New scanning and gene technology is allowing scientists to identify the disease at its earliest stages, often 15 years before symptoms appear and brain cells are destroyed, with drug trials in Colombia, USA and Europe showing startling success. The programme also reveals the changes in lifestyle that can prevent the development of the disease, as well as the effects of a UK-wide trial.
BBC2|1464046500|The Vikings Uncovered|||0|0|History|Dan Snow is joined by space archaeologist Dr Sarah Parcak to search for evidence of Viking settlements in North America, trying to prove that they settled in the New World 500 years before Columbus. Dan explores how they travelled west as first raiders, then settlers and traders throughout Britain and beyond to Iceland and Greenland, before excavating what could be the most westerly settlement ever discovered.(n)
BBC2|1464051900|Mary Beard's Ultimate Rome: Empire Without Limit|||1|3|Documentary|Scholar Mary Beard takes an in-depth look at identity and citizenship within the Roman Empire, including what it meant to be, or become, Roman, and how the different parts of the Empire reacted to Roman rule. She follows the story of an African Roman from his native land to Britain, where he served as a governor, and in York and Newcastle she finds the remains of Romans, but not as one might imagine.(n)
BBC2|1464055500|This Is BBC Two|||0|0|General Show,Game Show|Preview of upcoming programmes from BBC Two.(n)
BBC2|1464066000|Flog It! Trade Secrets|Tools of the Trade - Part One||2|3|Antiques,Collectibles|Paul Martin and the show's experts offer more advice on making money from antiques and collectibles, with this edition focusing on rare and valuable tools. There is also a feature on a piece of fascinating social history.(n)
BBC2|1464067800|Council House Crackdown|||2|1|General Education,Science|New series. The return of the programme that follows local authority housing officers as they track down social housing cheats, beginning with Croydon Council investigating a fraudulent tenant. Luke Doonan and Michelle Ackerley present.(n)
BBC2|1464070500|Family Finders|||0|0|General Education,Science|New series. The work of Britain's ever-growing army of commercial tracing companies and independent genealogy detective agencies. Together with more established bodies such as the Salvation Army, these dedicated staff devote their time to tracking down and reuniting lost family members.(n)
BBC2|1464073200|The Hairy Bikers' Pubs That Built Britain|Liverpool||1|6|Advertisement,Shopping|Si King and Dave Myers head to Liverpool, where they take a tour of some of the Swinging Sixties most important pubs. They meet John Lennon's drinking buddies from the 1950s to find out what he got up to over a pint or two before he was famous, discover why one pub was a regular for stars including Cilla Black, Gerry and the Pacemakers and the Beatles, and perform on stage at the Cavern Club.(n)
BBC2|1464075000|Great British Railway Journeys|Hampton Court to Teddington||7|19|General Education,Science|Michael Portillo starts his latest tour as Hampton Court Palace, where he is treated to a private tour of the Great Vine - the world's longest grapevine - before moving on to stately Claremont House, where tragic circumstances led directly to the birth of the Victorian era. He then moves up the line to Wimbledon and the site of a historic duelling event before ending his journey in Teddington, where he hears the story of a reformer whose work revolutionised the care for those with living disabilities.(n)
BBC2|1464076800|Victoria Derbyshire|24/05/2016||0|0|News Magazine,Current Affairs|Daily news and current-affairs programme offering discussion of breaking stories, exclusive interviews and audience interaction via social media.(n)
BBC2|1464084000|BBC Newsroom Live|24/05/2016||0|0|General News,Current Affairs|A chance to stay up to date on the day's leading stories, with the latest breaking news as it happens.(n)
BBC2|1464087600|Daily Politics|24/05/2016||0|0|Discussion,Debate|Parliamentary proceedings interspersed with discussions, interviews and filmed reports from around the country. Presented by Jo Coburn.(n)
BBC2|1464091200|The Super League Show|||0|0|Rugby League - Domestic|Tanya Arnold introduces action from the latest round of Super League matches, which saw every fixture take place at St James' Park in Newcastle on `Magic Weekend'.(n)
BBC2|1464093900|A Taste of Britain|Essex||1|5|Cooking|Janet Street-Porter and Brian Turner visit Mersea Island in Essex to learn about its culinary traditions and heritage. The pair chat to an oyster farmer whose family has been farming the same beds for decades and Brian cooks the shellfish for Janet to sample. He then meets fellow chef Darren Bennett at the Magic Mushroom where he serves up a meal of local trout before meeting pigs that produce prize-winning sausages. Meanwhile, Janet explores the history and geography of Cudmore Grove's unspoilt stretch of coastline.(n)
BBC2|1464096600|The TV That Made Me|Pam Ayres||1|11|Popular Culture,Traditional Arts|Brian Conley invites Pam Ayres to pick the TV shows that shaped her life, with the poet's selection including one of the scariest series ever broadcast on British TV.(n)
BBC2|1464098400|Holiday of My Lifetime with Len Goodman|Gloria Hunniford||1|12|Tourism,Travel|Gloria Hunniford revisits the town of Newcastle in Co Down to reminisce about a childhood holiday in 1948. She and presenter Len Goodman head to the hotel room she stayed in, walk in the Mourne Mountains and tuck into an Ulster fry-up and afternoon tea, before playing rounders on the beach.(n)
BBC2|1464101100|Caribbean with Simon Reeve|||1|1|Documentary|The adventurer travels around the islands and mainland coast of the Caribbean Sea, beginning on Hispaniola. He joins the Dominican Republic police's anti-narcotics division, before crossing the border to Haiti to see the notorious tented slums of Cite Soleil, while also discovering a vibrant, colourful and thriving side to the country. He ends this leg of his journey in Puerto Rico, an archipelago that is a territory of the United States, and examines the legacy of bombing and weapons testing on the island of Vieques.(n)
BBC2|1464104700|Great British Railway Journeys|Southport to Leyland||5|2|General Education,Science|Michael Portillo continues his journey around north-west England in the elegant resort town of Southport, where the railways provided thousands of holidaymakers with the chance enjoy the fun of the fair. On his journey around some of the region's larger towns, the presenter uncovers the history of Victorian entrepreneurship in Wigan and the beginnings of the Industrial Revolution in Bolton, before heading to smaller Leyland to get behind the wheel of a 100-year-old commercial vehicle.(n)
BBC2|1464106500|Bargain Hunt|Kedleston 29||36|14|Antiques,Collectibles|Antiques experts David Harper and Catherine Southon help two teams search for collectibles at a fair in the 820-acre parkland surrounding Kedleston Hall in Derbyshire. Meanwhile, Tim Wonnacott finds an unusual piece of Victoriana.(n)
BBC2|1464108900|Referendum Campaign Broadcast|Stronger IN Europe Campaign Broadcast||0|0|General Social,Political Issues,Economics|A referendum broadcast by the Stronger in Europe campaign, ahead of the Referendum on the United Kingdom's membership of the European Union, on June 23rd.(n)
BBC2|1464109200|Eggheads|||17|60|Game Show,Quiz|Jeremy Vine hosts the quiz in which the winners of famous game shows including Mastermind and Who Wants to Be a Millionaire? work as a team to tackle a new set of challengers hoping to win a cash prize.(n)
BBC2|1464111000|Countryfile Spring Diaries|A Sense of Spring!||1|2|Rural,Agricultural|Keeley Donovan discovers how just one in 50 people in the UK experiences Spring as a truly multi-sensory experience, and Margherita Taylor meets a man on a mission to make the countryside open to all.(n)
BBC2|1464112800|Antiques Road Trip|||12|0|Antiques,Collectibles|It's the final leg for Christina Trevanion and Thomas Plant. Kicking off from Gwersyllt in Wrexham, they meander through the border counties of Wales and England, buying antiques on their way. Their last auction takes place in Stoke-on-Trent, Staffordshire, before Charles Hanson and Margie Cooper embark on their trip from Melton Mowbray in Leicestershire to a Nottingham auction.(n)
BBC2|1464116400|RHS Chelsea Flower Show 2016|||1|6|Gardening|It's medals day at the RHS and Monty Don and Joe Swift reveal the show garden designs that have won a gold medal, as well as talking to the designer who has picked up the Best Show Garden award. Plus, news correspondent Kate Adie talks to Monty about her new-found passion for gardening.(n)
BBC2|1464120000|Old School with the Hairy Bikers|||1|3|Cooking|Si King and Dave Myers have four weeks left at the Oxford Academy to prove that their social experiment pairing up teenagers with pensioners is working. But there's trouble brewing. Jacub, who has ADHD, is still getting detentions and risks being thrown out of Old School unless he improves his behaviour. His older partner Clive is on a mission to find out how Jacub's gaming habit is affecting his learning. Last in the series.(n)
BBC2|1464123600|Later Live - with Jools Holland|||48|6|General Music,Ballet,Dance|The Last Shadow Puppets perform tracks from their recent chart-topping album Everything You've Come to Expect, while Californian singer-songwriter and slide guitar player Bonnie Raitt showcased her 20th album Dig in Deep. Plus, tracks by Malian kora player Ballake Sissoko and French cellist Vincent Segal, east London neo-soul singer Nao, veteran American alt-rock band Dinosaur Jr and Italian singer-songwriter Zucchero.(n)
BBC2|1464125400|Newsnight|24/05/2016||0|0|News Magazine,Current Affairs|Analysis of the day's events, presented by Emily Maitlis.(n)
BBC2|1464127800|Weather|||0|0|Weather|
BBC2|1464128100|Caravanner of the Year|||1|1|General|Six motorhome, caravan and camper van enthusiasts battle it out in the Caravan Club's inaugural competition to become Caravanner of the Year. Over two days, the contestants will take part in an awning assembly speed trial, before they are pushed to their limits by some challenging manoeuvres. Then, after competitive polishing and primping in the Concours D'Elegance, Chairman of the Caravan Club Grenville Chamberlain, journalist and motorhome maverick Andy Harris, and guest judge Lucy Jayne Grout choose the three who have earned a place in the final.(n)
BBC4|1463873400|Rod Stewart Live at Hyde Park|||0|0|General Music,Ballet,Dance|A concert by the singer that closed Radio 2's annual Festival in a Day, held in September 2015 in London's Hyde Park. Featuring a selection of hits from his back catalogue including Angel, In a Broken Dream, The Killing of Georgie (Part I and II) as well as Faces classics including Ooh La La and blues standard Rollin' and Tumblin'.
BBC4|1463877000|Top of the Pops: 1981|||0|0|Pop|Mike Read presents the October 1 edition, featuring music by the Tweets, Toyah, Altered Images, Gidea Park, the Creatures, Bad Manners, Dollar and Adam and the Ants.
BBC4|1463879400|Top of the Pops: 1981|||0|0|Pop|David `Kid' Jensen introduces an edition from October 1981, featuring performances by BA Robertson and Maggie Bell, the Exploited, Squeeze, Dave Stewart and Barbara Gaskin, This Year's Blonde, Toyah, Altered Images, Godley & Creme, the Creatures and Bad Manners. Plus, a dance sequence by Legs & Co.
BBC4|1463881800|Rod Stewart at the BBC|||0|0|General Music,Ballet,Dance|A tribute to the singer's career with a selection of his performances and interviews at the BBC. Songs include Sailing, You're in My Heart, I Don't Want to Talk About It and Da Ya Think I'm Sexy? Plus, Handbags and Gladrags from Rod's set at Glastonbury in 2002, his cover of Dorothy Fields' classic I'm in the Mood for Love and a song from his Radio 2 concert in May 2013.
BBC4|1463940000|Karajan's Magic and Myth|||0|0|General Education,Science|Documentary profiling Herbert von Karajan, arguably one of the most high-profile conductors in the history of classical music, exploring the many paradoxes in the life of this controversial figure. The Austrian was famed for his off-duty activities on the ski slopes, piloting his own jet, sailing his yacht, and driving fast cars, yet was a solitary man who enjoyed walking in the mountains. This programme examines his belief in the power of music, and his determination to leave behind a substantial legacy on film and features interviews with those who worked closely with him, including singers Placido Domingo and Jessye Norman, violinist Anne-Sophie Mutter, conductors Nikolaus Harnoncourt and Sir Neville Marriner, and the flautist Sir James Galway.
BBC4|1463945400|EastEnders|16/10/1986||0|0|Soap,Melodrama|A classic episode of the soap from 1986 directed by acclaimed film-maker Antonia Bird, which was the first episode of the show to feature only two characters. Den Watts has demanded a divorce from his wife Angie, who resorts to desperate measures to ensure he does not leave her. Starring Anita Dobson and Leslie Grantham.
BBC4|1463947200|From EastEnders to Hollywood: Antonia Bird|||0|0|Documentary|Profile of the director, whose career successful spanned the Royal Court Theatre, BBC dramas including Casualty and EastEnders to movies Safe, Priest, Face and Ravenous, before her death in 2013 at the age of 62. The programme explores the struggles she faced and the stories behind her movies, and features contributions from collaborators including Kay Mellor, Robert Carlyle, Anita Dobson and Irvine Welsh.
BBC4|1463952600|Care||2000|0|0|General Movie,Drama|A man struggles to piece together his life after suffering years of abuse in a children's home, a personal battle made doubly difficult by crusading reporters determined to expose the scandal. Drama directed by Antonia Bird and starring Steven Mackintosh, Jaye Griffiths and Charlotte Cornwell.
BBC4|1463958900|Horizon|Horizon: The Core||48|4|Documentary|Documentary following the scientists conducting experiments that try to recreate the conditions in Earth's core, an area 4,000 miles below the surface where storms rage in a sea of white-hot metal and a giant forest of crystals occupies a space the size of the moon.
BBC4|1463962500|Pop! The Science of Bubbles|||0|0|Documentary|Physicist Helen Czerski investigates the significance of bubbles, which can help to push back the boundaries of science, despite often being thought of as toys. She explores how a single one can reveal the workings of nature on a vast scale, and examines how globules of air formed as a result of breaking waves help oceans to breathe. The presenter also takes a look at the role bubbles are playing in the future design of ships and with new forms of medical treatment.
BBC4|1463966100|Karajan's Magic and Myth|||0|0|General Education,Science|Documentary profiling Herbert von Karajan, arguably one of the most high-profile conductors in the history of classical music, exploring the many paradoxes in the life of this controversial figure. The Austrian was famed for his off-duty activities on the ski slopes, piloting his own jet, sailing his yacht, and driving fast cars, yet was a solitary man who enjoyed walking in the mountains. This programme examines his belief in the power of music, and his determination to leave behind a substantial legacy on film and features interviews with those who worked closely with him, including singers Placido Domingo and Jessye Norman, violinist Anne-Sophie Mutter, conductors Nikolaus Harnoncourt and Sir Neville Marriner, and the flautist Sir James Galway.
BBC4|1464026400|World News Today|23/05/2016||0|0|News|The day's leading stories.
BBC4|1464028200|The Brecon Beacons with Iolo Williams|Winter||1|1|Nature,Animals|Iolo Williams explores the unique scenery of the Brecon Beacons over the course of a year, braving the elements in every season to detail the ever-changing landscape of the valleys. He begins in the winter, enduring a raging blizzard on the high peaks while the lowlands are bathed in sun. On the snowy slopes, foxes search for food while the great grey shrike - a ruthless hunter from Scandinavia - seeks other animals to eat. Plus, Iolo tracks red deer to the secluded gullies in one of the Beacons' wildest locations.
BBC4|1464030000|Dan Cruickshank: At Home with the British|The Cottage||1|1|Documentary|The historian celebrates British homes, starting with a visit to the picturesque Warwickshire countryside and the village of Stoneleigh, which has barely changed in 500 years, its cottages perfectly preserved. Here he charts the cottage's transformation from humble hovel to modern dream home.
BBC4|1464033600|Storm Troupers: The Fight to Forecast the Weather|||1|1|Documentary|New series. Journalist Alok Jha charts the history of weather forecasting from its origins in the early 19th century to the modern day, investigating how it was transformed from superstition into science. He reveals how pioneer Robert Fitzroy was driven by a desire to prevent disasters at sea, issuing Britain's first storm warnings and devising the first forecast to be published in a newspaper.
BBC4|1464037200|David Attenborough's Zoo Quest in Colour|||0|0|Nature,Animals|A one-off special showcasing colour footage from the 1950s wildlife series that launched the career of a young David Attenborough as a nature presenter. Using new-found film and behind-the-scenes stories from Attenborough and cameraman Charles Lague, this programme features clips of the best of Zoo Quest to West Africa, Zoo Quest to Guiana and Zoo Quest for a Dragon.
BBC4|1464042600|The Dark Ages: An Age of Light|The Men of the North||1|4|Documentary|In the final programme, Waldemar Januszczak turns his attention to the north of Europe, examining how Vikings marked their territory with rune stones, and decorated their long ships with intricate embellishment. He also investigates the jewellery and manuscript illumination created by the Irish and Anglo-Saxons, and examines how the Carolingians forecast their future as successors to Rome in the art they left behind. Last in the series.
BBC4|1464046200|Order and Disorder with Jim Al-Khalili|Information||1|2|General Education,Science|The theoretical physicist investigates the concept of information, exploring how humanity harnessed the power of symbols, including the first alphabet and the electric telegraph, through to the modern digital age. He also discovers how information is transmitted every day in many different forms, and is not solely reliant on human communication.(n)
BBC4|1464049800|Bullets, Boots and Bandages: How to Really Win at War|Stealing a March||1|2|History|Military historian Saul David explains the importance of efficiently moving an army during wartime, as he continues his exploration of the often-overlooked logistical issues that can make a major difference to the outcomes of conflicts. He also examines how generals have approached the problem in the past.(n)
BBC4|1464053400|The Brecon Beacons with Iolo Williams|Winter||1|1|Nature,Animals|Iolo Williams explores the unique scenery of the Brecon Beacons over the course of a year, braving the elements in every season to detail the ever-changing landscape of the valleys. He begins in the winter, enduring a raging blizzard on the high peaks while the lowlands are bathed in sun. On the snowy slopes, foxes search for food while the great grey shrike - a ruthless hunter from Scandinavia - seeks other animals to eat. Plus, Iolo tracks red deer to the secluded gullies in one of the Beacons' wildest locations.(n)
BBC4|1464055200|Storm Troupers: The Fight to Forecast the Weather|||1|1|Documentary|Journalist Alok Jha charts the history of weather forecasting from its origins in the early 19th century to the modern day, investigating how it was transformed from superstition into science. He reveals how pioneer Robert Fitzroy was driven by a desire to prevent disasters at sea, issuing Britain's first storm warnings and devising the first forecast to be published in a newspaper.(n)
BBC4|1464112800|World News Today|24/05/2016||0|0|News|The day's leading stories.(n)
BBC4|1464114600|The Brecon Beacons with Iolo Williams|Spring||1|2|Nature,Animals|Nesting season is in full swing as spring arrives and while hundreds of dotterel are resting in the Black Mountains during their journey from Africa to breeding sites in Scotland, peregrines are already nesting in an old quarry in the Central Beacons. Iolo Williams also explores the most crooked church in Britain and an old gunpowder works and finds that a 300-year-old stone wall reveals the history of this landscape.(n)
BBC4|1464116400|Storm Troupers: The Fight to Forecast the Weather|||1|1|Documentary|Journalist Alok Jha charts the history of weather forecasting from its origins in the early 19th century to the modern day, investigating how it was transformed from superstition into science. He reveals how pioneer Robert Fitzroy was driven by a desire to prevent disasters at sea, issuing Britain's first storm warnings and devising the first forecast to be published in a newspaper.(n)
BBC4|1464120000|Storyville|Last Days in Vietnam||0|0|Documentary|Oscar-nominated documentary about the final weeks of the Vietnam War, when the North Vietnamese Army closed in on Saigon as the panicked South Vietnamese people desperately attempted to escape. Including recollections of people who were there at the time.(n)
BBC4|1464125700|World War Two: 1945 & the Wheelchair President|||0|0|History|David Reynolds examines the wartime leadership of US president Franklin Roosevelt, who was burdened by secrets about his failing health and strained marriage.(n)
CBBC|1463896800|Arthur|The Pageant Pickle||18|19|Cartoons,Puppets|Arthur is excited when school ends for the summer, but first DW must have her Spring Pageant.
CBBC|1463897700|Scream Street|Mother of All Scares||1|5|General Children's,Youth|When Luke goes home to find that Otto has moved in, he must find out why he is there and how to get rid of him. He discovers Otto fled Sneer Hall to avoid a visiting relative with a temper, but when Luke brings her round so the two can reconcile, it does not quite go to plan.
CBBC|1463898300|Zig and Zag|DI Why?||1|2|Cartoons,Puppets|The alien twin brothers become DIY experts and set about fixing everything in Burb Street, regardless of whether it needs fixing or not.
CBBC|1463898900|Danger Mouse|Greenfinger||1|3|Cartoons,Puppets|Danger Mouse's attempts at gardening lead to a gigantic Welsh space plant taking over the world and an attack of intergalactic bees. Only Penfold's jam obsession can save the day!.
CBBC|1463899800|Dragons: Riders of Berk|What Flies Beneath||1|14|General Children's,Youth|Toothless tries to settle a score with an old rival, but Hiccup has to stop him before the encounter turns fatal. Children's entertainment spin-off series from the movie How to Train Your Dragon, following the adventures of Hiccup and his dragon.
CBBC|1463901000|Whoops I Missed the Bus|||3|8|General Children's,Youth|Revisiting CBBC's highlights from the past week, including Junior Vets on Call 2, Hetty Feather and Officially Amazing.
CBBC|1463902200|Ultimate Brain|Brain Factor!||2|5|General Children's,Youth|Science Super Hero Dr. Brain challenges three teams to prove that they have the Ultimate Brain. Finalists from X Factor 2014 - Stevi Ritchie, Betsy-Blue English and Parisa Tarjomani - take on two young teams in a mash up of science, entertainment and insanity. Today Guinea Pig tries to walk across some balancing beams while dodging a washing line, buckets and a giant fan - but has he got the S Factor?.
CBBC|1463904000|Blue Peter|||0|0|General Children's,Youth|The team presents a special edition allowing members of the BP fan club to control the show, with online votes, viewer comments and a chance to become Fans of the Month.
CBBC|1463905800|All Over the Workplace|Football||1|5|General Children's,Youth|Freya sees herself as a full-time professional footballer and Chitua wants to be a player before progressing to manager. They visit a professional football club where they are put through their paces by the coaches, then meet the manager to find out all about formations and tactics. Presented by Alex Riley.
CBBC|1463907600|Newsround|22/05/2016 - 1||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.
CBBC|1463907900|Matilda and the Ramsay Bunch|The Drive In||2|2|General Children's,Youth|The Cookie Monster pays a surprise visit, so Matilda Ramsay gets his help and together they set to work making a giant chocolate-chip treat. The Ramsay Bunch has planned a drive-in movie night in the back garden, and as darkness falls its members set to work. Along with their friend Cruz Beckham they build the outdoor screen, while Matilda cooks margherita and pepperoni pizza with a rainbow salad. As well as cooking, Matilda makes a prank film and the whole family falls for her tricks - even dad Gordon.
CBBC|1463908800|The Next Step|Don't Stop the Party||2|1|General Children's,Youth|The A-Troupe is reunited after their win at regionals, while Emily and Michelle set aside their differences over Eldon.
CBBC|1463910300|Lost & Found Music Studios|Day After Day||1|7|Drama|John is having trouble at home and decides to move into the band's van, much to Luke's dismay. Clara gets stage fright when she tries to perform with other members of the studio.
CBBC|1463911800|Our School|In Trouble||1|4|General Children's,Youth|Year seven student Ewan's behaviour challenges his teachers at his new school.
CBBC|1463913600|The Dengineers|Hawaiian Den||1|4|General Children's,Youth|Mark Wright and Lauren Layfield come to the aid of Ella, who would love a Hawaiian-style beach hut getaway to help her escape a family home filled with 35 bikes.
CBBC|1463915400|Newsround|22//05/2016 - 2||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.
CBBC|1463915700|All Over the Place: USA|||1|4|Entertainment - Teens|Ed Petrie, Iain Stirling, Richard Whisker, Naomi Wilkinson, Barney Harwood, Ceallach Spellman and Michelle Ackerley set out to find the most unusual, strange and amazing places to visit in the United States of America. They ride a rollercoaster that is housed inside the country's largest shopping mall, cross seven miles of ocean on one of the world's longest bridges, and embark on a road trip to a classic car and bike museum.
CBBC|1463917500|Horrible Histories|||5|6|Comedy|Queen Victoria's coronation fails to go according to plan, George IV takes part in Historical Come Dine with Me, and Alexander the Great refuses to stop conquering things.
CBBC|1463919000|Marrying Mum and Dad|1980s||2|9|General Children's,Youth|Naomi Wilkinson and Ed Petrie help Cassie and Marnie plan a 1980s-themed Jewish wedding for their mum and stepdad, who get to drive a DeLorean - made famous in Back to the Future.
CBBC|1463920800|Naomi's Nightmares of Nature|South Africa: North||1|2|Nature,Animals|Naomi Wilkinson tracks down dangerous fauna living in the savannahs of northern South Africa, and goes in search of one of the biggest creatures on Earth.
CBBC|1463922600|Newsround|22/05/2016 - 3||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.
CBBC|1463922900|4 O'Clock Club|Time Capsule||4|7|Comedy|Nero and the gang decide to sabotage parents' evening, while Josh finds out the truth about his missing dad.
CBBC|1463924700|How to Be Epic @ Everything|||1|2|Entertainment - Teens|Children's series in which experts show how they do their specialist skills, including playing rock guitar, spinning a basketball, grooming a horse and skimming a stone.
CBBC|1463925600|Hank Zipzer|Ballot Box Blunder||2|7|Comedy|When a seat on the school council becomes available, Hank uses charm, personality and his mum's pastries to try to stop it from going to McKelty. However, Emily attempts to win the election another way - by convincing everybody that she's too cool for school.
CBBC|1463927100|Hank Zipzer|Valentine's Confusion||2|8|Comedy|Hank has his heart set on asking Anya to the Valentine's dance, but soon discovers that this year Valentine's Day is doing funny things to people and he ends up in a pickle when he tries to please more than one girl. Meanwhile, Rosa and Stan are proving that even as grown-ups Valentine's can be a confusing time - if only there were rules?.
CBBC|1463928600|Hank Zipzer|Camouflage||2|9|Comedy|With Emily in hospital having her tonsils out and a history project due, Hank decides the best possible course of action is to take Katherine - Emily's lizard and best friend - into school. Meanwhile at the hospital, Stan is trying to prove to Rosa that he's not squeamish - easier said than done when all you want to do is pass out.
CBBC|1463930100|Hank Zipzer|Hank's Birthday||2|10|Comedy|It's Hank's 13th birthday and he wants the greatest party of all time. Unfortunately Stan and Rosa have other ideas, so Hank decides to have a secret party of his own in the den. Nothing can go wrong with that - right?.
CBBC|1463931600|Hank Zipzer|Hank's New School||2|11|Comedy|After yet another bad parents' evening, Stan is determined to get Hank a good education - at another school. Desperate not to leave Frankie, Ashley and Mr Rock behind, Hank is forced to do the unthinkable and fight to stay at Westbrook Academy. Mr Rock, on the other hand, finds an old friend's offer of a life away from Westbrook extremely tempting.
CBBC|1463933100|Hank Zipzer|Papa Pete In Love||2|12|Comedy|When Hank gets a B-plus at school thanks to even more of Papa Pete's support he realises he owes his grandad big time and gets the idea to find him a new girlfriend. What could go wrong? Back at home, Emily has a new boyfriend and a suspicious Stan grills him about his intentions he realises his mistake.
CBBC|1463934900|Hank Zipzer|Last Day||2|13|Comedy|Hank is determined to make it through the last day of term without a detention - but an incident with an egg in assembly changes all of that and he finds himself in danger of being excluded from school permanently. Comedy, starring Nick James and Henry Winkler.
CBBC|1463936400|The Dengineers|Hawaiian Den||1|4|General Children's,Youth|Mark Wright and Lauren Layfield come to the aid of Ella, who would love a Hawaiian-style beach hut getaway to help her escape a family home filled with 35 bikes.
CBBC|1463938200|Copycats|||4|2|Games and Quizzes|Alfie's team from the Vale of Glamorgan go up against Liani's team from East London, battling it out for a chance to get to the Ballroom and play for the Copycats trophy. Game show, presented by Sam Nixon and Mark Rhodes.
CBBC|1463940000|Hetty Feather|Strike||1|6|Drama|Nurse Winston is sacked by Matron so Hetty convinces the children to go on strike.
CBBC|1463941800|Eve|Things That Go Beep in the Night||1|6|Drama|Eve goes to a Halloween party and makes a friend in good-looking Zac. Nick discovers that Katherine has found a way to track down the location of the military chip inside Eve placing Project Eternity in jeopardy, so tries to throw her off the scent.
CBBC|1463943600|Deadly 60|Mexico 1||3|6|General Children's,Youth|Steve Backshall chases sailfish in Mexico's Yucatan Peninsula, and dives on a pristine reef in search of a real-life sea monster.
CBBC|1463945400|Junior Bake Off|||1|6|Cooking|The cooks race to bake a lemon drizzle cake in one hour and create a recipe based on the theme of America. Meanwhile, Aaron Craze finds out about cupcakes.
CBBC|1463983200|Arthur|Some Assembly Required||18|20|Cartoons,Puppets|DW cannot wait to test out her new play set, but she has to settle for just the box and her imagination while the toy is being built.
CBBC|1463983800|Sidekick|Ice to Know You||1|31|General Children's,Youth|Eric turns summer into winter and threatens to start a new ice age.
CBBC|1463984700|Danger Mouse|The Unusual Suspects||1|13|Cartoons,Puppets|When secret information is leaked from HQ all eyes fall on Colonel K! Is it possible he's a traitor or is there something suspicious about him moustache?.
CBBC|1463985600|Newsround|23/05/2016 - 1||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.
CBBC|1463985900|Officially Amazing|||5|6|Entertainment - Pre-Teens|The Moffat brothers return and hope to break yet another motoring record. Presented by Ben Shires, Haruka Kuroda and Al Jackson.
CBBC|1463986800|How to Be Epic @ Everything|||1|7|Entertainment - Teens|Experts show how to perform a skateboard trick, shuffle cards, make a shelter and survive being bitten by a venomous snake.
CBBC|1463987700|Newsround|23/05/2016 - 2||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.
CBBC|1463988300|Tracy Beaker Returns|Big Brother||3|4|General Children's,Youth|Liam is tagged for a crime he did not commit, then a letter arrives from someone claiming to be his long lost brother. Comedy based on the books by Jacqueline Wilson.
CBBC|1463990100|Hank Zipzer|Battle of the Goblins||1|4|Comedy|The accident-prone boy breaks his and Frankie's science project, and then messes up when trying to collect a game for his friend. He finally thinks he may have finally found a solution to his problems - but disaster strikes again.
CBBC|1463991600|Help! My Mini School Trip Is Magic|The Broomstick||1|4|General Children's,Youth|John is clearing up at the dogs' home when his assistant unexpectedly ends up flying high on a broomstick.
CBBC|1463991900|Roy|Pint-Sized Roy||2|6|Cartoons,Puppets|The cartoon boy is accidentally shrunk and destroys the anniversary cake Becky baked for their grandparents.
CBBC|1463993700|Naomi's Nightmares of Nature|Yucatan||3|8|Nature,Animals|Naomi Wilkinson explores Mexico's Yucatan peninsula, where she plays Russian roulette, meets a master of disguise, and witnesses a spectacle of nature - an army of over two million bats.
CBBC|1463995500|Ice Stars|The Big Decision||1|2|General Children's,Youth|Josh is struggling to land his jumps, and speed skater Maddie has a new plan as she attempts to recover from a mystery illness.
CBBC|1463997000|Marrying Mum and Dad|Army||4|2|General Children's,Youth|A tank is the wedding transport and an assault course is the entertainment for this surprise army-themed wedding. Hosted by Naomi Wilkinson and Ed Petrie.
CBBC|1463998800|Wolfblood|Morwal||4|4|General Children's,Youth|Jana's uneasy relationship with Imara is tested during a mission to find a dangerous wolfblood. Supernatural drama, starring Leona Vaughan.
CBBC|1464000600|The Next Step|Winner Takes It All||1|30|General Children's,Youth|The team goes up against Elite Studios at the final of the regional competition, and Michelle and Eldon work hard to perfect their duo.
CBBC|1464001800|Hank Zipzer|Battle of the Goblins||1|4|Comedy|The accident-prone boy breaks his and Frankie's science project, and then messes up when trying to collect a game for his friend. He finally thinks he may have finally found a solution to his problems - but disaster strikes again.
CBBC|1464003600|Ice Stars|The Big Decision||1|2|General Children's,Youth|Josh is struggling to land his jumps, and speed skater Maddie has a new plan as she attempts to recover from a mystery illness.
CBBC|1464005100|Naomi's Nightmares of Nature|Yucatan||3|8|Nature,Animals|Naomi Wilkinson explores Mexico's Yucatan peninsula, where she plays Russian roulette, meets a master of disguise, and witnesses a spectacle of nature - an army of over two million bats.
CBBC|1464006900|Marrying Mum and Dad|Army||4|2|General Children's,Youth|A tank is the wedding transport and an assault course is the entertainment for this surprise army-themed wedding. Hosted by Naomi Wilkinson and Ed Petrie.
CBBC|1464008700|Tracy Beaker Returns|Big Brother||3|4|General Children's,Youth|Liam is tagged for a crime he did not commit, then a letter arrives from someone claiming to be his long lost brother. Comedy based on the books by Jacqueline Wilson.
CBBC|1464010500|Officially Amazing|||5|6|Entertainment - Pre-Teens|The Moffat brothers return and hope to break yet another motoring record. Presented by Ben Shires, Haruka Kuroda and Al Jackson.
CBBC|1464011400|How to Be Epic @ Everything|||1|7|Entertainment - Teens|Experts show how to perform a skateboard trick, shuffle cards, make a shelter and survive being bitten by a venomous snake.
CBBC|1464012300|Shaun the Sheep|Big Top Timmy||1|16|Cartoons,Puppets|A circus sets up in a nearby field, and a spellbound Timmy wanders off to investigate. Can Shaun rescue him before the farmer notices he's gone?.
CBBC|1464012600|Shaun the Sheep|Fetching||1|17|Cartoons,Puppets|Bitzer falls in love with a female from the local camp-site, but the flock creates havoc in the farmhouse, forcing Shaun to get the sheepdog's mind back on his job.
CBBC|1464013200|Sidekick|Maxum Man Mark 2||1|1|General Children's,Youth|The adventures of four students at the Academy for Aspiring Sidekicks. In the first episode, Eric and Trevor try to clone Maxum Man, but inadvertently create a creature that is half-human, half-hamster.
CBBC|1464013800|OOglies|||1|1|Cartoons,Puppets|Lonely Sprout looks for a vegetable friend, and the see-sawing grapes try to avoid an invasion by clumsy Melonhead.
CBBC|1464014700|Zig and Zag|School Rules||1|5|Cartoons,Puppets|The alien brothers go to school to learn how to solve a crossword clue, causing classroom chaos all the way to the bell.
CBBC|1464015600|Just Kidding|||1|26|Comedy|Children's comedy show that lets them concoct pranks to play on unsuspecting adults.
CBBC|1464016800|Newsround|23/05/2016 - 3||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.
CBBC|1464017400|Lost & Found Music Studios|Sunrise||1|12|Drama|Maggie's uncle offers the girls a chance to open for one of their favourite bands, but there's a big catch, while Clara is having trouble dealing with the aftermath of the plagiarism scandal. Isaac is disappointed to learn that his brother, underground hip-hop producer Tully, is dating Mary and spending more time at Lost & Found.
CBBC|1464018900|Lifebabble|Cyberbullying||1|7|General Children's,Youth|The team tackles cyberbullying, revealing how easy it is to unintentionally victimise people online. Chavala and Dr Aaron are also on hand to offer advice and guidance to viewers.
CBBC|1464019200|All Over the Workplace|Police||1|7|General Children's,Youth|Alex Riley follows the fortunes of Abi and Kyra as the tackle the world of law enforcement, apprehending a car thief and arresting a bank robber.
CBBC|1464021000|The Dumping Ground|Holding On||2|6|Drama|Expectations are high when Tyler's mum pays a visit. Drama based on books by Jacqueline Wilson, starring Connor Byrne and Kay Purcell.
CBBC|1464022800|Zig and Zag|Meet the Robo-Parents||1|6|Cartoons,Puppets|The duo create Robo-parents simply to use them to get the family deal at the Pizzeria. However, the robots' parental programme gets out of control.
CBBC|1464023400|Endangered Species|Merl's Birthday Curse||1|32|Cartoons,Puppets|When Merl is convinced his birthday is cursed because he has never had a good birthday party, Pickle and Gull try to make this year's party the best ever.
CBBC|1464024300|Dragons: Riders of Berk|In Dragons We Trust||1|5|General Children's,Youth|The dragons are blamed for a crime outbreak, so Hiccup sets out to discover what is really going on before they are exiled.
CBBC|1464025500|Danger Mouse|Sinistermouse||2|3|Cartoons,Puppets|When an evil version of Danger Mouse escapes from a parallel dimension and joins forces with Baron Greenback, the hero may have finally met his match.
CBBC|1464026400|Horrible Histories|||3|5|Comedy|Louis XVI and Marie Antoinette go on Historical Wife Swap with some French peasants, and Queen Cleopatra sings about her femme fatale reputation. A Welsh prince from the Middle Ages endures a very stupid death and a Tudor peasant gets a makeover in Historical Fashion Fix.
CBBC|1464028200|Operation Ouch|||4|2|General Children's,Youth|The doctors reveal where blood comes from, Dr Chris meets a patient undergoing life-changing brain surgery, and there's a mind-bending trick to test the powers of concentration. There are also more medical mysteries in 'Ouch & About', and in Accident & Emergency one patient's in with a double sporting injury while another has taken a nasty tumble with her horse.
CBBC|1464030000|Epic Quick Blast|||2|5|Entertainment - Pre-Teens|How to make giant smoke rings, harmonise and pull off a cool football trick.
CBBC|1464030300|The Next Step|Winner Takes It All||1|30|General Children's,Youth|The team goes up against Elite Studios at the final of the regional competition, and Michelle and Eldon work hard to perfect their duo.
CBBC|1464031800|The Dumping Ground|Mischief||3|4|Drama|Bailey finally finds a friend while battling to adopt a homeless dog. Drama based on books by Jacqueline Wilson, starring Connor Byrne and Kay Purcell.(n)
CBBC|1464069600|Arthur|Shelter from the Storm - Part One||19|1|Cartoons,Puppets|Part one of two. A hurricane hits Elwood City and everyone is affected. Ladonna's father is called up by the army corps of engineers, while Arthur struggles to reunite lost pets and owners.(n)
CBBC|1464070200|Sidekick|Graduation Daze||1|99|General Children's,Youth|The aspiring heroes finally graduate from the Academy for Aspiring Sidekicks.(n)
CBBC|1464071100|Danger Mouse|Danger Fan||1|14|Cartoons,Puppets|A visit of the crimebusting rodent's biggest fan coincides with members of the team starting to disappear. Revival of the classic cartoon, with the voice of Alexander Armstrong.(n)
CBBC|1464072000|Newsround|24/05/2016 - 1||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.(n)
CBBC|1464072300|Officially Amazing|||5|7|Entertainment - Pre-Teens|Gymnast and stuntman Alex Jerram attempts a twisting vault record.(n)
CBBC|1464073200|How to Be Epic @ Everything|||1|8|Entertainment - Teens|Experts reveal how to do sign language, make ice-cream, launch a rocket and handle a crab. Narrated by Cel Spellman.(n)
CBBC|1464074100|Newsround|24/05/2016 - 2||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.(n)
CBBC|1464074700|Tracy Beaker Returns|Belonging||3|5|General Children's,Youth|Tracy gets tangled up in Lily's plan to reunite Poppy and Rosie with their dad. Meanwhile, a stray three-legged dog attaches itself to Frank.(n)
CBBC|1464076500|Hank Zipzer|Haunted Hank||1|5|Comedy|Emily is picked on by Nick McKelty, prompting Hank to seek revenge by building the world's scariest haunted house in a bid to give the bully the fright of his life.(n)
CBBC|1464078000|Help! My Mini School Trip Is Magic|The Ballerina||1|5|General Children's,Youth|In this episode, twinkle-toed trickster Katherine is at the Royal Opera House.(n)
CBBC|1464078300|Roy|A Crushing Blow||2|7|Cartoons,Puppets|The cartoon boy wonders whether he could be falling in love with Kathy, his arch nemesis.(n)
CBBC|1464080100|Naomi's Nightmares of Nature|Bonus Bits||3|9|Nature,Animals|Naomi Wilkinson shares unseen bonus highlights from the filming of series three, including the lethal leap of the biggest big cat in Finland, searching the spooky jungles of Borneo for a toxic teddy and a colony of giant bats in Thailand.(n)
CBBC|1464081900|Ice Stars|The Sin Bin||1|3|General Children's,Youth|Ice hockey teammates Liam and Rais have the biggest match of the season. While Rais is doing some training with his dad, Liam is determined to keep a lid on his combative style.(n)
CBBC|1464083400|Marrying Mum and Dad|Prehistoric||4|3|General Children's,Youth|Elle and her friends plan a prank-filled prehistoric wedding where the couple exchange their vows in a cave while dressed as cavemen.(n)
CBBC|1464085200|Wolfblood|The Quiet Hero||4|5|General Children's,Youth|TJ tries to help Selina with a problem that threatens to expose her as a wolfblood. Starring Rukku Nahar.(n)
CBBC|1464087000|The Next Step|Don't Stop the Party||2|1|General Children's,Youth|The A-Troupe is reunited after their win at regionals, while Emily and Michelle set aside their differences over Eldon.(n)
CBBC|1464088200|Hank Zipzer|Haunted Hank||1|5|Comedy|Emily is picked on by Nick McKelty, prompting Hank to seek revenge by building the world's scariest haunted house in a bid to give the bully the fright of his life.(n)
CBBC|1464090000|Ice Stars|The Sin Bin||1|3|General Children's,Youth|Ice hockey teammates Liam and Rais have the biggest match of the season. While Rais is doing some training with his dad, Liam is determined to keep a lid on his combative style.(n)
CBBC|1464091500|Naomi's Nightmares of Nature|Bonus Bits||3|9|Nature,Animals|Naomi Wilkinson shares unseen bonus highlights from the filming of series three, including the lethal leap of the biggest big cat in Finland, searching the spooky jungles of Borneo for a toxic teddy and a colony of giant bats in Thailand.(n)
CBBC|1464093300|Marrying Mum and Dad|Prehistoric||4|3|General Children's,Youth|Elle and her friends plan a prank-filled prehistoric wedding where the couple exchange their vows in a cave while dressed as cavemen.(n)
CBBC|1464095100|Tracy Beaker Returns|Belonging||3|5|General Children's,Youth|Tracy gets tangled up in Lily's plan to reunite Poppy and Rosie with their dad. Meanwhile, a stray three-legged dog attaches itself to Frank.(n)
CBBC|1464096900|Officially Amazing|||5|7|Entertainment - Pre-Teens|Gymnast and stuntman Alex Jerram attempts a twisting vault record.(n)
CBBC|1464097800|How to Be Epic @ Everything|||1|8|Entertainment - Teens|Experts reveal how to do sign language, make ice-cream, launch a rocket and handle a crab. Narrated by Cel Spellman.(n)
CBBC|1464098700|Shaun the Sheep|Mountains out of Molehills||1|18|Cartoons,Puppets|A freshly dug molehill spoils the flock's fun, and Shaun has to resort to extreme measures to get rid of the pesky mole.(n)
CBBC|1464099000|Shaun the Sheep|Buzz Off Bees||1|13|Cartoons,Puppets|The sheep discover a mysterious buzzing object in their field - so Shaun investigates and finds it is full of bees.(n)
CBBC|1464099600|Sidekick|To Party Perchance to Party||1|2|General Children's,Youth|Eric and Trevor try to crash Vana's party while fighting the villian Drilliam Shakespeare.(n)
CBBC|1464100200|OOglies|||1|2|Cartoons,Puppets|The soaps indulge their love of extreme sports as they make their way to the living room, and Mr Magnetic attracts trouble in the form of mischievous tinfoil.(n)
CBBC|1464101100|Zig and Zag|Meet the Robo-Parents||1|6|Cartoons,Puppets|The duo create Robo-parents simply to use them to get the family deal at the Pizzeria. However, the robots' parental programme gets out of control.(n)
CBBC|1464102000|Just Kidding|||2|1|Comedy|Children's comedy show that lets them concoct pranks to play on unsuspecting adults.(n)
CBBC|1464103200|Newsround|24/05/2016 - 3||0|0|General Children's,Youth|Current affairs reports aimed at a younger audience.(n)
CBBC|1464103800|Hetty Feather|Words from Home||2|3|Drama|Hetty has a surprise visitor with important news.(n)
CBBC|1464105600|Marrying Mum and Dad|Jungle||1|5|General Children's,Youth|Ed Petrie and Naomi Wilkinson help two boys organise a jungle-themed wedding for their parents, complete with lemurs and lions.(n)
CBBC|1464107400|The Dumping Ground|Endurance||2|7|Drama|A very long night ensues when two opposing Dumping Ground teams take up a bizarre telly challenge. Drama based on books by Jacqueline Wilson, starring Connor Byrne and Kay Purcell.(n)
CBBC|1464109200|Zig and Zag|Fanzillas||1|7|Cartoons,Puppets|The alien twin brothers become football superfans, but they learn that it is all about the winning, and not just the taking part, as they cost Burbia United the cup.(n)
CBBC|1464109800|Endangered Species|Speechless||1|33|Cartoons,Puppets|Merl finds a switch that turns off Pickle's voice. He loves the peace and quiet at first, but soon misses his pals' playful racket.(n)
CBBC|1464110700|Dragons: Riders of Berk|Alvin and the Outcasts||1|6|General Children's,Youth|Alvin and the outcast Vikings terrorise Berk, which has been left defenceless without its dragons. Hiccup is the only one who can bring them back.(n)
CBBC|1464111900|Danger Mouse|There's No Place Like Greenback||1|20|Cartoons,Puppets|DM and Penfold become reluctant parents when it appears the Baron has wiped his own memory. With the voices of Alexander Armstrong and Kevin Eldon.(n)
CBBC|1464112800|Horrible Histories|||3|6|Comedy|Henry VIII demonstrates his diet of all meat and no vegetables, and Bob Hale tries to explain the War of the Roses, which took place in the Middle Ages. Plus, a Stone Age man invents farming, and Admiral Nelson causes confusion with his last words.(n)
CBBC|1464114600|Operation Ouch|||4|3|General Children's,Youth|With the help of opera singer Lucy O'Bryne, the Doctors reveal the hidden muscle that makes you breathe, Dr Xand heads to a DNA laboratory to solve the mystery of who stole his strawberry milk, and there's a chance to play along at home with another mind-bending trick. Meanwhile, the 'Ouch Mobile' is open for business, and over in Accident & Emergency one patient has cut their eyebrow, and another has stapled his own finger.(n)
CBBC|1464116400|Epic Quick Blast|||2|6|Entertainment - Pre-Teens|Tips on how to become a gymnast, fold a T-shirt in one second, and cook snails.(n)
CBBC|1464116700|The Next Step|Don't Stop the Party||2|1|General Children's,Youth|The A-Troupe is reunited after their win at regionals, while Emily and Michelle set aside their differences over Eldon.(n)
CBeebies|1463893200|Show Me Show Me|Scarecrows and Statues||5|3|General Children's,Youth|Chris, Pui and all the other toys explore the outside world, and Miss Mouse finds a helpful scarecrow to look after her crops.
CBeebies|1463894400|Justin's House|House for Sale||2|6|General Children's,Youth|Robert and Little Monster concoct a plan to stop Justin selling his house.
CBeebies|1463895900|Baby Jake|Baby Jake Loves Bouncing Apples||1|14|General Children's,Youth|Nibbles the rabbit joins Jake in the orchard, and the friends have fun bouncing.
CBeebies|1463896800|Raa Raa the Noisy Lion|Ooo Ooo's Wriggly Jiggly Game||2|8|General Children's,Youth|The cub organises a series of games for Topsy's party, but not everybody is good at them.
CBeebies|1463897400|Postman Pat: SDS|Postman Pat and the Chinese Dragon||2|14|General Children's,Youth|Pumpkin scares the locals by getting his head stuck in a Chinese dragon costume, and it is up to Pat to calm everyone down and deliver the outfit to school in time for Chinese Day.
CBeebies|1463898300|Dinopaws|The Thing That Fell Down||1|5|Cartoons,Puppets|Bob wishes to see one of the twinkles in the night sky up close. Animated adventures with the three young dinosaurs Bob, Gwen and Tony.
CBeebies|1463898900|Hey Duggee|The Paper Boat Badge||1|16|Cartoons,Puppets|The dog's newspaper boat blows away and the squirrels race to rescue it.
CBeebies|1463899200|Chuggington|Wilson and the Ice-Cream||1|25|General Children's,Youth|Wilson is asked to take refrigerated cars to the ice-cream fair, but when Frostini offers him a tour of the factory, he forgets about his important job.
CBeebies|1463899800|Octonauts|Yeti Crab||3|8|Cartoons,Puppets|Tweak tests the Gup-X down in the midnight zone, but a yeti crab damages the ship putting both itself and the octonauts in danger.
CBeebies|1463900700|Kate & Mim-Mim|Super Kate||1|41|Cartoons,Puppets|Kate wonders what it is like to have superpowers when she gets her ball stuck in a tree, while in Mimiloo, Tack reveals a new supercharger invention and Boomer is in a predicament.
CBeebies|1463901300|Everything's Rosie|Will at the Wheel||4|15|General Children's,Youth|Will converts his old potters wheel to make Holly a present.
CBeebies|1463901900|Peter Rabbit|The Tale of the Mystery Plum Thief||1|16|General Children's,Youth|It appears that a thief has beaten Peter to the last plum on Mr McGregor's tree.
CBeebies|1463902800|Tree Fu Tom|The Great Journey||1|16|General Children's,Youth|Tom and Twigs get a crash course in being Ranchers and have to lead a baby beetle drive on their own.
CBeebies|1463904000|Something Special|Something Special: Out and About: Zookeeper||7|20|General Children's,Youth|Justin and his friends help out at the zoo, and Mr Tumble discovers what it is like to be an animal.
CBeebies|1463905200|Chuggington: Badge Quest|Chug Patrol||1|4|General Children's,Youth|The friends try to break the record for the number of problems reported on the rails, as they go on a chug patrol to earn another badge.
CBeebies|1463905500|Our Family|Meet Raphael and Eli's Family||1|14|General Children's,Youth|Meet brothers, 5-year old Raphael and 3-year old Eli. They love vegetables, so decide to visit a neighbour's allotment to pick their own. But who's going to fix the broken wheelbarrow? And what will they find amongst the worms? At home, they make something very special with the beetroot they have brought back from the allotment - beetroot chocolate brownies! So 'chefs', Raphael and Eli get down to some baking!.
CBeebies|1463906400|Footy Pups|Penalties||1|14|General Children's,Youth|Arsenal player Rachel Yankey and her team take part in a gripping penalty shootout. Meanwhile, Rozzie struggles to score against a team of stinky Skunks. Narrated by John Motson.
CBeebies|1463907300|Topsy and Tim|Big Box||1|11|General Children's,Youth|The duo cannot wait to find out what is inside the box that they have taken care of for Mr Fishwick.
CBeebies|1463907900|Topsy and Tim|Finders Seekers||1|12|General Children's,Youth|The twins play hide-and-seek with their friends, but Rai becomes stuck in the bathroom.
CBeebies|1463908500|Jamillah and Aladdin|The Eggless Chicken||1|6|General Children's,Youth|Aladdin is heartbroken when his mother orders him to take his favourite chicken, Warqa to the butcher's shop. However, Jamillah has a plan, and with Genie's help they find a way to make Warqa the most valuable chicken of all.
CBeebies|1463909400|Octonauts|The Swashbuckling Swordfish||2|14|Cartoons,Puppets|Kwazii explores a pirate shipwreck that is guarded by three swashbuckling swordfish while searching for a mythical sword.
CBeebies|1463910300|Peter Rabbit|The Tale of the Hazelnut Raid||1|23|General Children's,Youth|Peter accidentally destroys the squirrels' store of nuts, and sets off to Owl Island to replace them.
CBeebies|1463910900|Spot Bots Zoople Time|The Musical Mermaids: Seaweedophone||1|14|Games and Quizzes|Laugh and play along with the Spot Bots with a quick game to get you switched on. Bubbles & Rock play some sounds on their funny Seaweedophone. Try to remember the right order of the sounds they play.
CBeebies|1463911200|Swashbuckle|The Daringly Dangerous Expedition||1|4|Games and Quizzes|Four youngsters aim to retrieve Gem's jewels and make one of the pirates walk the plank. Meanwhile, Cook and Line's manage to ruin Captain Stinker's plans for a grand adventure.
CBeebies|1463912700|Gigglebiz|||2|8|General Children's,Youth|Singing waiter Opera Oliver plays `gooseberry' between two romantic diners, King Flannel helps the butler to wash the royal car and Gail Force presents a world transport exclusive from Little Bottom station. Live-action comedy sketch show for the under-sixes, starring Justin Fletcher.
CBeebies|1463913600|Mister Maker's Arty Party|||1|15|Pre-School|How to make fabulous furry monster pictures, and how artist Salvador Dali painted monster-like creatures in his works of art.
CBeebies|1463914800|Melody|Storm||2|14|General Children's,Youth|Mum and Melody visit Shoreham Lifeboat Station. Mum says she has some music for Melody to listen to called Storm Interlude from Peter Grimes, by Benjamin Britten.
CBeebies|1463915400|Balamory|I Spy||1|63|Pre-School|The children on Edie's bus get bored, but Josie Jump and PC Plum are on hand to entertain them.
CBeebies|1463916600|I Can Cook|Frittata||1|23|General Children's,Youth|The children visit the garden to learn how asparagus grows, before cooking Italian frittatas. Presented by Katy Ashworth.
CBeebies|1463917500|Grandpa in My Pocket|A Saturday Full of Surprises||1|22|Comedy|Grandpa tries to make a grumpy Great Aunt Loretta laugh when she comes round and spoils his plans for a Saturday afternoon playing with Jason.
CBeebies|1463918400|My Story|Polo||2|16|General Children's,Youth|A man shares his memories with his daughter, including his life growing up in Kenya and his love of horses and playing polo. Narrated by Nicky Campbell.
CBeebies|1463919300|Tilly and Friends|Flighty-Bitey||1|16|General Children's,Youth|Doodle spoils a picnic in the garden when he eats too much cake.
CBeebies|1463919900|Waybuloo|Whizzcrackers||1|24|Pre-School|Yoyojo keeps missing the whizzcrackers that appear in the sky, so everyone makes whizzybongles by throwing bongleberries up in the air.
CBeebies|1463921100|Big Barn Farm|Hide & Seek||1|16|Cartoons,Puppets|The farmyard gang plays a game of hide and seek.
CBeebies|1463922000|Something Special|Something Special: Out and About: Zookeeper||7|20|General Children's,Youth|Justin and his friends help out at the zoo, and Mr Tumble discovers what it is like to be an animal.
CBeebies|1463923200|Chuggington: Badge Quest|Chug Patrol||1|4|General Children's,Youth|The friends try to break the record for the number of problems reported on the rails, as they go on a chug patrol to earn another badge.
CBeebies|1463923500|Our Family|Meet Raphael and Eli's Family||1|14|General Children's,Youth|Meet brothers, 5-year old Raphael and 3-year old Eli. They love vegetables, so decide to visit a neighbour's allotment to pick their own. But who's going to fix the broken wheelbarrow? And what will they find amongst the worms? At home, they make something very special with the beetroot they have brought back from the allotment - beetroot chocolate brownies! So 'chefs', Raphael and Eli get down to some baking!.
CBeebies|1463924400|Footy Pups|Penalties||1|14|General Children's,Youth|Arsenal player Rachel Yankey and her team take part in a gripping penalty shootout. Meanwhile, Rozzie struggles to score against a team of stinky Skunks. Narrated by John Motson.
CBeebies|1463925300|Topsy and Tim|Big Box||1|11|General Children's,Youth|The duo cannot wait to find out what is inside the box that they have taken care of for Mr Fishwick.
CBeebies|1463925900|Topsy and Tim|Finders Seekers||1|12|General Children's,Youth|The twins play hide-and-seek with their friends, but Rai becomes stuck in the bathroom.
CBeebies|1463926500|Jamillah and Aladdin|The Eggless Chicken||1|6|General Children's,Youth|Aladdin is heartbroken when his mother orders him to take his favourite chicken, Warqa to the butcher's shop. However, Jamillah has a plan, and with Genie's help they find a way to make Warqa the most valuable chicken of all.
CBeebies|1463927400|Octonauts|The Swashbuckling Swordfish||2|14|Cartoons,Puppets|Kwazii explores a pirate shipwreck that is guarded by three swashbuckling swordfish while searching for a mythical sword.
CBeebies|1463928000|Peter Rabbit|The Tale of the Hazelnut Raid||1|23|General Children's,Youth|Peter accidentally destroys the squirrels' store of nuts, and sets off to Owl Island to replace them.
CBeebies|1463928900|Spot Bots Zoople Time|The Musical Mermaids: Seaweedophone||1|14|Games and Quizzes|Laugh and play along with the Spot Bots with a quick game to get you switched on. Bubbles & Rock play some sounds on their funny Seaweedophone. Try to remember the right order of the sounds they play.
CBeebies|1463929200|Justin's House|The Wishing Wardrobe||1|20|General Children's,Youth|Justin is very excited to discover a fancy dress day is taking place in Justin Town, and wonders what to wear.
CBeebies|1463930700|Andy's Wild Adventures|Cheetahs||2|20|General Children's,Youth|Andy and Kip embark on a wild adventure to Africa in search of the world's fastest land mammal - the cheetah.
CBeebies|1463931600|Mister Maker's Arty Party|||1|15|Pre-School|How to make fabulous furry monster pictures, and how artist Salvador Dali painted monster-like creatures in his works of art.
CBeebies|1463932800|Swashbuckle|The Daringly Dangerous Expedition||1|4|Games and Quizzes|Four youngsters aim to retrieve Gem's jewels and make one of the pirates walk the plank. Meanwhile, Cook and Line's manage to ruin Captain Stinker's plans for a grand adventure.
CBeebies|1463934300|Sarah & Duck|Slow Quest||1|27|Cartoons,Puppets|Tortoise embarks a mission through Sarah and Duck's house, so the pair try to work out what he is crawling toward.
CBeebies|1463934600|Katie Morag|Katie Morag and the Carrot Competition||2|5|General Children's,Youth|Neilly Beag and Grannie Island hold a competition to see who can grow the biggest carrot, but the challenge brings unexpected results.
CBeebies|1463935500|Katie Morag|Katie Morag and the Big Shinty Match||2|6|General Children's,Youth|Struay must win their upcoming shinty match against Coll to keep the cup, so Neilly Beag trains extra hard to make sure he is picked for the team.
CBeebies|1463936400|Clangers|Space Tangle||1|11|Cartoons,Puppets|Small notices that the Iron Chicken has become trapped by junk metal that has got caught in orbit around her nest, but Major comes up with a clever solution.
CBeebies|1463937000|The Adventures of Abney & Teal|Rock Music||2|26|General Children's,Youth|The duo must find a way to compromise when Abney is trying to write poetry, but Teal just wants to make noise.
CBeebies|1463937600|In the Night Garden|Upsy Daisy, Igglepiggle, the Bed and the Ball||1|29|Cartoons,Puppets|Igglepiggle decides to sleep in Upsy Daisy's bed while she plays with a ball in the garden.
CBeebies|1463939400|CBeebies Bedtime Story|Chocolate Mousse - Nadia Hussain||0|0|Pre-School|Nadia Hussain reads Chocolate Mousse for Greedy Goose, by Julia Donaldson.
CBeebies|1463979600|Show Me Show Me|Trombones and Jumpers||5|4|General Children's,Youth|The Tiddlers help Mr Bloom make a cloche to keep his pepper seedlings warm, while inside the nursery Sebastian has received a postcard from his mother.
CBeebies|1463980800|Justin's House|Back in Time||2|7|General Children's,Youth|Justin entertains children with singing, dancing and comedy, assisted by Robert the robot butler, Little Monster and unicycling delivery lady, Dee Livery.
CBeebies|1463982300|Raa Raa the Noisy Lion|Wake Up Huffty||2|19|General Children's,Youth|Huffty fails to appear as the other animals gather to listen to the dawn chorus, so Raa Raa and his friends try to wake him so he can enjoy the event.
CBeebies|1463983200|Teletubbies|Taking a Ride||1|41|Pre-School|The friends ride the Dup Dup and the Tubby Custard Machine also takes them for a jaunt. In Tummy Tales, a boy goes on a cable car.
CBeebies|1463984100|Bing|Toy Party||2|40|Cartoons,Puppets|The bunny gets jealous when Sula gives Pando more attention on a playdate. He tries to gain some for himself and ends up being pushed, so Amma show them how to get rid of the anger.
CBeebies|1463984700|Hey Duggee|The Cake Badge||1|2|Cartoons,Puppets|Happy decides to eat a cake they have found in a field, but they are unsure who its real owner is.
CBeebies|1463985000|Boj|Gavin's Got Talent||1|36|Cartoons,Puppets|The friends put on a talent show, but Gavin's act the Mega-Robot-Dancer 64i does not work and the event cannot continue - so Boj tries to persuade him he has his own special talent.
CBeebies|1463985600|The Furchester Hotel|Toast with a Smile||1|7|General Children's,Youth|Elmo must deliver a tray of toast to a hungry guest, but along the way must dodge the horses, trolleys, bumps in the rug and monsters.
CBeebies|1463986500|Octonauts|The Dwarf Lanternshark||1|44|Cartoons,Puppets|Captain Barnacles and the team try to find an injured dwarf lanternshark.
CBeebies|1463987100|Mike the Knight|Viking Snow Day||1|51|Cartoons,Puppets|The youngster discovers that Vikings have landed in Glendragon and is sure they have come to cause trouble.
CBeebies|1463988000|Charlie and Lola|I Can't Stop Hiccupping||3|10|Cartoons,Puppets|Lola's concert preparations are interrupted when she gets the hiccups.
CBeebies|1463988600|Rastamouse|Da Cool Cruiser||1|10|Cartoons,Puppets|The Easy Crew investigates when a mischievous mouse breaks Zoomer's skates and steals wheels from Fats' garage.
CBeebies|1463989200|Nelly & Nora|Cold in the Bed||1|10|General Children's,Youth|Nelly suffers a bout of sickness and is confined to bed, so Nora tries to cheer her up. Animation about the adventures of two sisters at a seaside camping park.
CBeebies|1463989800|Mr Bloom: Here and There|Down to Earth Farm||2|16|Cartoons,Puppets|Mr Bloom meets Drew and Felicia who show him how to milk a goat, collect eggs from chickens and harvest tomatoes and sweetcorn. Plus, they make a scarecrow for the vegetable garden.
CBeebies|1463990400|My First|Potty||1|17|General Children's,Youth|In this episode we follow Ellis as she starts potty training.
CBeebies|1463991000|Bing|Skateboard||2|17|Cartoons,Puppets|Flop and Bing visit the park where they see Pando on a skateboard and decide to try it out for themselves - but discover that it is much harder to balance than it looks.
CBeebies|1463991600|Bing|Toy Party||2|40|Cartoons,Puppets|The bunny gets jealous when Sula gives Pando more attention on a playdate. He tries to gain some for himself and ends up being pushed, so Amma show them how to get rid of the anger.
CBeebies|1463991900|Wussywat the Clumsy Cat|Heavy||1|32|Cartoons,Puppets|The curious cat discovers the difference between heavy and light objects when he helps Ortus stop his seed packets from blowing away.
CBeebies|1463992500|Twirlywoos|Pulling||2|30|Pre-School|Great BigHoo, Toodloo, Chickedy and Chick have a tug-of-war with a carpenter when they pull on the end of her tape measure. Back in the Boat, the Twirlywoos find a vine coming out of Peekaboo's house, and cannot resist giving it a pull.
CBeebies|1463993100|Something Special|Something Special: We're All Friends: Shopping||9|23|General Children's,Youth|Justin and his friends go on a bus trip to the shops, and Mr Tumble sets up his own outlet at home.
CBeebies|1463994300|Let's Play|Ancient Roman||2|5|Education|Rebecca discovers whether she has what it takes to be an ancient Roman as she helps builders Cementicus and Fabulous finish the Emperor's new villa.
CBeebies|1463995500|Mister Maker Around the World|||1|23|General Children's,Youth|There is an attempt to make an apple surprise against the clock, while in South America, the Mini Makers build a crocodile swamp, and get inspiration from a giraffe in South Africa.
CBeebies|1463996700|Ruff-Ruff, Tweet and Dave|A Rainbow Adventure||1|23|General Children's,Youth|The trio learn all the colours of the rainbow by naming and matching colours in Hatty's garden.
CBeebies|1463997300|Tinga Tinga Tales|Why Caterpillar Is Never in a Hurry||1|9|Cartoons,Puppets|Animals rush around to get ready for a parade, while Caterpillar is happy to sit in a tree and munch on leaves.
CBeebies|1463998200|Magic Hands|Daffodils||2|6|General Children's,Youth|A mysterious flute leads Donna and Ashley on a musical adventure in which Pink Bird dresses up as Pan to play sweet tunes and all the creatures dress up as daffodils.
CBeebies|1463998800|My Pet and Me|Goldfish||2|11|General Children's,Youth|Rory helps Thomas change the water in his goldfish's tank and they also give the pet some food.
CBeebies|1463999700|Minibeast Adventure with Jess|Moth||1|16|General Children's,Youth|Zoologist Jess French learns about moths, and sets up a trap overnight in a bid to collect some of the more beautiful varieties.
CBeebies|1464000000|Waybuloo|A Surprise for Yojojo||2|2|Pre-School|Yojojo's drum skin breaks, so his fellow Piplings decide to surprise him by fixing it and decorating his bandstand.
CBeebies|1464001200|Melody|Who's at the Door?||2|16|General Children's,Youth|Mum takes Melody to visit a cathedral. The partially sighted girl feels the carved wooden door, picking out different shapes. She asks Mum for some church door music, and Beethoven's Symphony No 5 is duly chosen.
CBeebies|1464001800|Balamory|Beach Ball||1|3|Pre-School|Josie wants to go to the beach, but first she has to overcome a minor problem.
CBeebies|1464003000|I Can Cook|Chunky Banana Bread||1|24|General Children's,Youth|Katy Ashworth is joined by junior cooks to find out how sugar is made and have fun making chunky banana bread.
CBeebies|1464003900|Grandpa in My Pocket|There Came a Big Spider||4|9|Comedy|Grandpa and Elsie make space spiders for their Captain Dumbletwit puppet play, but it all proves too much for Great Aunt Loretta.
CBeebies|1464004800|My First|Potty||1|17|General Children's,Youth|In this episode we follow Ellis as she starts potty training.
CBeebies|1464005400|Bing|Skateboard||2|17|Cartoons,Puppets|Flop and Bing visit the park where they see Pando on a skateboard and decide to try it out for themselves - but discover that it is much harder to balance than it looks.
CBeebies|1464006000|Bing|Toy Party||2|40|Cartoons,Puppets|The bunny gets jealous when Sula gives Pando more attention on a playdate. He tries to gain some for himself and ends up being pushed, so Amma show them how to get rid of the anger.
CBeebies|1464006300|Wussywat the Clumsy Cat|Heavy||1|32|Cartoons,Puppets|The curious cat discovers the difference between heavy and light objects when he helps Ortus stop his seed packets from blowing away.
CBeebies|1464006900|Twirlywoos|Pulling||2|30|Pre-School|Great BigHoo, Toodloo, Chickedy and Chick have a tug-of-war with a carpenter when they pull on the end of her tape measure. Back in the Boat, the Twirlywoos find a vine coming out of Peekaboo's house, and cannot resist giving it a pull.
CBeebies|1464007500|Something Special|Something Special: We're All Friends: Shopping||9|23|General Children's,Youth|Justin and his friends go on a bus trip to the shops, and Mr Tumble sets up his own outlet at home.
CBeebies|1464008700|Let's Play|Ancient Roman||2|5|Education|Rebecca discovers whether she has what it takes to be an ancient Roman as she helps builders Cementicus and Fabulous finish the Emperor's new villa.
CBeebies|1464009900|Mister Maker Around the World|||1|23|General Children's,Youth|There is an attempt to make an apple surprise against the clock, while in South America, the Mini Makers build a crocodile swamp, and get inspiration from a giraffe in South Africa.
CBeebies|1464011100|Ruff-Ruff, Tweet and Dave|A Rainbow Adventure||1|23|General Children's,Youth|The trio learn all the colours of the rainbow by naming and matching colours in Hatty's garden.
CBeebies|1464011700|Tinga Tinga Tales|Why Caterpillar Is Never in a Hurry||1|9|Cartoons,Puppets|Animals rush around to get ready for a parade, while Caterpillar is happy to sit in a tree and munch on leaves.
CBeebies|1464012600|Magic Hands|Daffodils||2|6|General Children's,Youth|A mysterious flute leads Donna and Ashley on a musical adventure in which Pink Bird dresses up as Pan to play sweet tunes and all the creatures dress up as daffodils.
CBeebies|1464013200|Tilly and Friends|Tumpty's Skipping Rope||1|45|General Children's,Youth|The pals play with hula hoops and go skipping, but Tumpty cannot fit through even the biggest hoop.
CBeebies|1464013800|Timmy Time|Timmy's Picnic||1|11|General Children's,Youth|The class enjoys a picnic and game of football, but when Apricot's spikes cause the ball to burst, she makes up for it by using them to pick up litter.
CBeebies|1464014400|Spot Bots|Zipperoo||1|10|Cartoons,Puppets|Get switched on and play games with the Spot Bots. Cubi is showing off with his rocket powered zip wire.
CBeebies|1464015600|Swashbuckle|The Big Fall Out||3|11|Games and Quizzes|Join Gem's daring Swashbucklers as they attempt to win back her jewels from the naughty pirates Cook, Line and Captain Sinker, in this hilarious and fast-paced physical gameshow. Cook and Line have fallen out so Captain Sinker needs to play the peace-maker and restore order. Meanwhile, Hermione, Maaria, Harrison and Josh are the Swashbucklers aiming to win back all Gem's jewels and earn the right to see one of the pirates walk the plank into the Ship's Mess!.
CBeebies|1464016800|Messy Goes to Okido|A Sock Too Far||1|42|Cartoons,Puppets|The monster and his friends go camping with a robot who can do anything.
CBeebies|1464017400|Andy's Prehistoric Adventures|Sabre-Toothed Cat & Roar||1|11|General Children's,Youth|Andy leaps into his time-traveling clock to visit a fearsome sabre-toothed cat, but when his gizmo malfunctions he is accidentally shrunk down to the size of an insect.
CBeebies|1464018300|Peter Rabbit|The Tale of the Tunnel Rumbler||2|5|General Children's,Youth|The rabbit and friends believe there is a mysterious invader in their tunnels, but getting rid of it proves to be difficult with Tommy Brock nearby.
CBeebies|1464019200|Tree Fu Tom|It's a Kind of Magic||3|4|General Children's,Youth|A red magic lesson goes badly wrong when Twigs breaks Muru's magic stick.
CBeebies|1464020700|Our Family|Noah Throws a Party for Sketch||2|9|General Children's,Youth|Four-year-old Noah throws a birthday party for his dog Sketch, hanging decorations and baking a cake with his dad, and making a card and wrapping a special present with his mum.
CBeebies|1464021300|Gigglebiz|||3|5|General Children's,Youth|Will Singalot infuriates the gang with his non-stop singing and Robin tries some log-walking to impress Maid Marion.
CBeebies|1464022200|Sarah & Duck|World Bread Day||1|28|Cartoons,Puppets|The youngster and her feathered friend take part in a treasure hunt when there is a bread festival in the park.
CBeebies|1464022800|Clangers|The Ball||1|29|Cartoons,Puppets|Tiny and Small find a strange silver ball that glows and rings when it bounces. Mother tells them it is a living thing, and Granny is convinced it must have friends nearby.
CBeebies|1464023400|The Adventures of Abney & Teal|The Porridge Party||1|1|General Children's,Youth|The duo make lots of porridge to warm themselves up on a cold and gloomy day, but soon realise they have produced too much.
CBeebies|1464024000|In the Night Garden|Tombliboo Ooo Drinks Everybody Else's Pinky Ponk Juice||1|30|Cartoons,Puppets|Tombliboo Ooo makes himself ill by drinking too much Pinky Ponk juice, so his friends play music to make him feel better.
CBeebies|1464025800|CBeebies Bedtime Story|When the Dragons Came - Aaron McCusker||0|0|Pre-School|Aaron McCusker reads When the Dragons Came, by Naomi Kefford and Lynne Moore.(n)
CBeebies|1464066000|Show Me Show Me|Confetti and Roadsweepers||5|5|General Children's,Youth|Chris and Pui cannot stop throwing confetti, and when there is far too much to sweep up, Miss Mouse comes to the rescue.(n)
CBeebies|1464067200|Justin's House|Posh Nosh||2|8|General Children's,Youth|Roberta the superturbo robot must try to fix Justin's Cake-a-pulter Hundred Thousand after Robert fails to do so, but not before Justin treats the duo to a not-so-peaceful dinner.(n)
CBeebies|1464068700|Raa Raa the Noisy Lion|The Lion's Share||2|20|General Children's,Youth|The animals try to work out what the new toy Raa Raa has made does.(n)
CBeebies|1464069600|Teletubbies|Photos||1|42|Pre-School|The friends take selfies with the Tubby Phone and a child in Tummy Tales has their photo taken in a photo booth with their grandparent.(n)
CBeebies|1464070500|Bing|Mobile Phone||2|38|Cartoons,Puppets|Bing is playing the talking lettuce game on Flop's phone when he drops the phone and accidentally breaks it. Too panicked to tell Flop what's he's done Bing puts the phone in the bin but he's so upset that Flop knows something has happened.(n)
CBeebies|1464071100|Hey Duggee|The Hair Badge||1|3|Cartoons,Puppets|Duggee is having a bad hair day, and the Squirrels may not be able to help him.(n)
CBeebies|1464071400|Boj|The Giggly Park Express||1|37|Cartoons,Puppets|The friends make a train for Denzil and his teddies using cardboard boxes, and go on a trip around the world.(n)
CBeebies|1464072000|The Furchester Hotel|Isabel Gets the Ding-Ups||1|8|General Children's,Youth|Isabel suffers from bell-monster hiccups and the Furchesters need to stop them so she can welcome all the guests with a friendly ding.(n)
CBeebies|1464072900|Octonauts|The Pirate Parrotfish||1|45|Cartoons,Puppets|The crew goes on a pirate treasure hunt and Kwazii meets the perfect sidekick - a parrotfish.(n)
CBeebies|1464073500|Mike the Knight|Mike the Knight and the Night Time Lookout||2|1|Cartoons,Puppets|Mike learns that even knights require naps when he falls asleep while serving as a lookout.(n)
CBeebies|1464074400|Charlie and Lola|But I Am Completely Hearing and Also Listening||3|11|Cartoons,Puppets|Lola resolves to learn to listen after her inattention gets her into trouble both at home and at school.(n)
CBeebies|1464075000|Rastamouse|Da Monstrous Fib||1|11|Cartoons,Puppets|The orphan mice are spooked by scary sounds during a camping trip, so Rastamouse has to reassure everyone that there are no such things as monsters.(n)
CBeebies|1464075600|Nelly & Nora|Blown Away||1|11|General Children's,Youth|It is too windy for umbrellas and hats, but not for Nelly and Nora.(n)
CBeebies|1464076200|Mr Bloom: Here and There|Hythe Ferry||2|17|Cartoons,Puppets|Mr Bloom meets three children who love the Hythe Ferry, and goes for a ride on an electric train. Together they draw a picture to be made into a plaque for a pier.(n)
CBeebies|1464076800|My First|Musical Experience||1|18|General Children's,Youth|Following Levi as he explores all of the songs and sounds in the world around him, and learns all about music, eventually finding his own favourite instrument.(n)
CBeebies|1464077400|Bing|Butterfly||2|18|Cartoons,Puppets|The bunny tries to help a butterfly that has flown inside the nursery and landed on Sula's painting.(n)
CBeebies|1464078000|Bing|Mobile Phone||2|38|Cartoons,Puppets|Bing is playing the talking lettuce game on Flop's phone when he drops the phone and accidentally breaks it. Too panicked to tell Flop what's he's done Bing puts the phone in the bin but he's so upset that Flop knows something has happened.(n)
CBeebies|1464078300|Wussywat the Clumsy Cat|Compost||1|33|Cartoons,Puppets|The feline helps Ortus plant his cabbages but they run out of compost. It remains to be seen where they will find some more.(n)
CBeebies|1464078900|Twirlywoos|Full||1|1|Pre-School|The friends eat too much and feel full, and after seeing someone pour water into a glass, they get carried away finding their own containers to fill.(n)
CBeebies|1464079500|Something Special|Something Special: We're All Friends: Cookery||9|24|General Children's,Youth|Justin and his friends prepare pizzas, while Mr Tumble wants to make a carrot cake.(n)
CBeebies|1464080700|Let's Play|Nurse||2|6|Education|Sid steps through the magic curtain and plays being a nurse. He must try to manage to look after a busy ward of sick patients and deal with a special visitor's injury.(n)
CBeebies|1464081900|Mister Maker Around the World|||1|24|General Children's,Youth|An attempt to make a card tube creature in less than a minute in Australia, while in the UK the Mini Makers help to create a mountain of cakes.(n)
CBeebies|1464083100|Ruff-Ruff, Tweet and Dave|An Exploring Adventure||1|24|General Children's,Youth|Ruff-Ruff, Tweet and Dave go exploring, following clues which lead them to discover a strange new animal - a `doggy-birdy-panda' that is a mixture of all three of them put together.(n)
CBeebies|1464083700|Tinga Tinga Tales|Why Mosquito Buzzes||1|10|Cartoons,Puppets|An African fable explaining why mosquitos make a buzzing sound when they fly.(n)
CBeebies|1464084600|Magic Hands|The Fairies||2|7|General Children's,Youth|Sheba the Snake and Click Clack the Crab take centre stage as Ashley and Aimee explore where fairies and elves live and what they do.(n)
CBeebies|1464085200|My Pet and Me|Ducks||2|12|General Children's,Youth|Ferne Corrigan visits Aaron and his pet ducks, and together they clean out their home and fill up the duck pond.(n)
CBeebies|1464086100|Minibeast Adventure with Jess|Spider||1|17|General Children's,Youth|Zoologist Jess French takes a look at some spiders, then accompanies a group of children to have a look for webs and eggs.(n)
CBeebies|1464086400|Waybuloo|Cheebie Tune||2|3|Pre-School|NokTok makes a music box, but does not think the last note sounds right, so all the Piplings help him look for a new piece of wood.(n)
CBeebies|1464087600|Melody|Music Box||2|17|General Children's,Youth|Mum and Melody discover Granny's broken music box, and Mum gives her Clair De Lune by Debussy, which captures the youngster's imagination.(n)
CBeebies|1464088200|Balamory|The Missing Scarecrow||1|4|Pre-School|PC Plum asks the children in the nursery to help him make a scarecrow.(n)
CBeebies|1464089400|I Can Cook|Katy's Lasagne||1|25|General Children's,Youth|Katy Ashworth and the team find out how mozzarella cheese is made, before using it to prepare a lasagne.(n)
CBeebies|1464090300|Grandpa in My Pocket|The Wonderbubble Weather Watcher||4|10|Comedy|Mr Mentor's new invention, The Wonderbubble Weather Watcher, reads that it is the perfect weather for a boat trip - but Grandpa is not so sure.(n)
CBeebies|1464091200|My First|Musical Experience||1|18|General Children's,Youth|Following Levi as he explores all of the songs and sounds in the world around him, and learns all about music, eventually finding his own favourite instrument.(n)
CBeebies|1464091800|Bing|Butterfly||2|18|Cartoons,Puppets|The bunny tries to help a butterfly that has flown inside the nursery and landed on Sula's painting.(n)
CBeebies|1464092400|Bing|Mobile Phone||2|38|Cartoons,Puppets|Bing is playing the talking lettuce game on Flop's phone when he drops the phone and accidentally breaks it. Too panicked to tell Flop what's he's done Bing puts the phone in the bin but he's so upset that Flop knows something has happened.(n)
CBeebies|1464092700|Wussywat the Clumsy Cat|Compost||1|33|Cartoons,Puppets|The feline helps Ortus plant his cabbages but they run out of compost. It remains to be seen where they will find some more.(n)
CBeebies|1464093300|Twirlywoos|Full||1|1|Pre-School|The friends eat too much and feel full, and after seeing someone pour water into a glass, they get carried away finding their own containers to fill.(n)
CBeebies|1464093900|Something Special|Something Special: We're All Friends: Cookery||9|24|General Children's,Youth|Justin and his friends prepare pizzas, while Mr Tumble wants to make a carrot cake.(n)
CBeebies|1464095100|Let's Play|Nurse||2|6|Education|Sid steps through the magic curtain and plays being a nurse. He must try to manage to look after a busy ward of sick patients and deal with a special visitor's injury.(n)
CBeebies|1464096300|Mister Maker Around the World|||1|24|General Children's,Youth|An attempt to make a card tube creature in less than a minute in Australia, while in the UK the Mini Makers help to create a mountain of cakes.(n)
CBeebies|1464097500|Ruff-Ruff, Tweet and Dave|An Exploring Adventure||1|24|General Children's,Youth|Ruff-Ruff, Tweet and Dave go exploring, following clues which lead them to discover a strange new animal - a `doggy-birdy-panda' that is a mixture of all three of them put together.(n)
CBeebies|1464098100|Tinga Tinga Tales|Why Mosquito Buzzes||1|10|Cartoons,Puppets|An African fable explaining why mosquitos make a buzzing sound when they fly.(n)
CBeebies|1464099000|Magic Hands|The Fairies||2|7|General Children's,Youth|Sheba the Snake and Click Clack the Crab take centre stage as Ashley and Aimee explore where fairies and elves live and what they do.(n)
CBeebies|1464099600|Tilly and Friends|The Five Tillys||1|46|General Children's,Youth|The friends imitate Tilly, but then start to miss being themselves.(n)
CBeebies|1464100200|Timmy Time|Timmy Tries to Hide||1|12|General Children's,Youth|Noisy Paxton ruins a game of hide-and-seek, so Timmy teaches him how to play, only to conceal himself so well the class cannot find him in time for snacks.(n)
CBeebies|1464100800|Spot Bots|Ziptastic Tower||1|11|Cartoons,Puppets|Cubi and Lexi try to build a perfect, but delicate, tower of bricks, and they cannot resist fiddling with their creation.(n)
CBeebies|1464102000|Swashbuckle|Plant Hunters||3|13|Games and Quizzes|Gem's team try to win back her jewels, while Captain Sinker challenges Cook and Line to find her a brand new flower so she can be like the plant-hunters of old.(n)
CBeebies|1464103200|Messy Goes to Okido|Rumbly Tummy||1|43|Cartoons,Puppets|Messy's tummy is rumbling and so is Lofty the giant's. Luckily the gang are hungry to solve this scientific mystery.(n)
CBeebies|1464103800|Andy's Prehistoric Adventures|Centrosaurus & Video||1|12|General Children's,Youth|Andy heads back in time to search a prehistoric forest for a plant-munching dinosaur, but runs into a relative of the T-rex instead, and then joins a herd of centrosaurus.(n)
CBeebies|1464104700|Peter Rabbit|The Tale of the Best Bowler||2|6|General Children's,Youth|A pine cone bowling rivalry between Peter and Nutkin gets out of hand and causes trouble.(n)
CBeebies|1464105600|Go Jetters|Table Mountain, South Africa||1|17|General Children's,Youth|Glitch wants to ski, so the Grimbots give Table Mountain a snowy peak, which threatens its rare plants.(n)
CBeebies|1464106200|Go Jetters|The Statue of Liberty, USA||1|7|General Children's,Youth|Grandmaster Glitch makes the Statue of Liberty fall, right into the path of a passing ferry.(n)
CBeebies|1464107100|Our Family|Charlotte and Zoe's Tea Party||2|12|General Children's,Youth|Sisters six-year old Charlotte and five-year old Zoe prepare a banana cake with Mum's help, then they invite Mum, Dad and their toys to a tea party to taste what they have made.(n)
CBeebies|1464107700|Gigglebiz|||3|6|General Children's,Youth|Incompetent DIY Dan demonstrates how to liven up a front door, gardener Will Barrow has trouble with a worm while trying to eat lunch, and antiques expert Ann Teak examines a rare pearl necklace.(n)
CBeebies|1464108600|Sarah & Duck|Pond Princess||1|29|Cartoons,Puppets|The ducks award Sarah a crown at the pond so she tries to work out what her royal duties should be.(n)
CBeebies|1464109200|Clangers|Planty||1|30|Cartoons,Puppets|The friends help Granny make her knitting space more special. Major makes her a fan and Mother gives her a purple plant from her garden called Planty. Michael Palin narrates.(n)
CBeebies|1464109800|The Adventures of Abney & Teal|Firefly Lullaby||1|6|General Children's,Youth|The Poc-Pocs keep waking Abney and Teal up during the night, and Neep encounters fireflies.(n)
CBeebies|1464110400|In the Night Garden|Looking for Each Other||1|31|Cartoons,Puppets|Igglepiggle cannot find Upsy Daisy and asks Makka Pakka for help.(n)
BBC News|1463871600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463873400|Reporters|||0|0|reserved|A weekly showcase of the best reports from the BBC's global network of correspondents.
BBC News|1463875200|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463877000|The Travel Show|21/05/2016||0|0|reserved|Join the team on their journey of discovery as they explore new destinations around the globe and uncover hidden sides to some of the world's favourite holiday hotspots.
BBC News|1463878800|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463880600|Dateline London|21/05/2016||0|0|reserved|Foreign correspondents currently posted to London look at events in the UK through outsiders' eyes, and at how the issues of the week are being tackled around the world.
BBC News|1463882400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463884200|Our World|21/05/2016||0|0|General Social,Political Issues,Economics|Global current affairs.
BBC News|1463886000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463887800|Click|21/05/2016||0|0|Computers,Internet,Gaming|A guide to the latest gadgets, websites, games and computer industry news.
BBC News|1463889600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463891400|The Week in Parliament|20/05/2016||0|0|General News,Current Affairs|A round-up of the week's proceedings in Parliament, presented by Alicia McCarthy.
BBC News|1463893200|Breakfast|||0|0|General Social,Political Issues,Economics|A round-up of national and international news, plus sports reports, weather forecasts and arts and entertainment features.
BBC News|1463896800|Breakfast|||0|0|News|Early-morning reports.
BBC News|1463900400|Breakfast|||0|0|News|Early-morning reports.
BBC News|1463904000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463905800|The Papers|22/05/2016 - 1||0|0|reserved|No need to wait until tomorrow morning to see what's in the papers - tune in to BBC News and hear a lively, informed and engaging conversation about the next day's papers.
BBC News|1463907600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463909400|Horizon|||0|0|Documentary|Series examining topical scientific issues.
BBC News|1463911200|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463913000|Dateline London|21/05/2016||0|0|reserved|Foreign correspondents currently posted to London look at events in the UK through outsiders' eyes, and at how the issues of the week are being tackled around the world.
BBC News|1463914800|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463916600|Click|21/05/2016||0|0|Computers,Internet,Gaming|A guide to the latest gadgets, websites, games and computer industry news.
BBC News|1463918400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463920200|The Travel Show|21/05/2016||0|0|reserved|Join the team on their journey of discovery as they explore new destinations around the globe and uncover hidden sides to some of the world's favourite holiday hotspots.
BBC News|1463922000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463923800|The Week in Parliament|20/05/2016||0|0|General News,Current Affairs|A round-up of the week's proceedings in Parliament, presented by Alicia McCarthy.
BBC News|1463925600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463927400|Click|21/05/2016||0|0|Computers,Internet,Gaming|A guide to the latest gadgets, websites, games and computer industry news.
BBC News|1463929200|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463931000|Talking Movies|||0|0|General Arts,Culture|News and reviews from the US cinema scene, with Tom Brook.
BBC News|1463932800|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463936400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463940000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463941800|Sportsday|||0|0|General Sports|Results and analysis from countrywide events.
BBC News|1463942700|Meet The Author|||0|0|reserved|Writers talk about their latest books.
BBC News|1463943600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463945400|The Travel Show|21/05/2016||0|0|reserved|Join the team on their journey of discovery as they explore new destinations around the globe and uncover hidden sides to some of the world's favourite holiday hotspots.
BBC News|1463947200|World News Today|22/05/2016||0|0|News|The day's leading stories.
BBC News|1463949000|Our World|21/05/2016||0|0|General Social,Political Issues,Economics|Global current affairs.
BBC News|1463950800|BBC News|22/05/2016||0|0|News|The latest national and international stories as they break.
BBC News|1463953500|The Papers|22/05/2016 - 2||0|0|reserved|No need to wait until tomorrow morning to see what's in the papers - tune in to BBC News and hear a lively, informed and engaging conversation about the next day's papers.
BBC News|1463954400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463956200|The Papers|22/05/2016 - 3||0|0|reserved|No need to wait until tomorrow morning to see what's in the papers - tune in to BBC News and hear a lively, informed and engaging conversation about the next day's papers.
BBC News|1463957100|The Film Review|20/05/2016||0|0|reserved|Mark Kermode gives his unique take on the best and worst of the week's film and DVD releases, with Gavin Esler.
BBC News|1463958000|Newsday|||0|0|News Magazine,Current Affairs|
BBC News|1463959800|Reporters|21/05/2016||0|0|reserved|A weekly showcase of the best reports from the BBC's global network of correspondents.
BBC News|1463961600|Newsday|||0|0|News Magazine,Current Affairs|
BBC News|1463963400|Asia Business Report|||0|0|News Magazine,Current Affairs|Live from Singapore the essential business news as it breaks and a look ahead to the news that will shape the business day.
BBC News|1463964300|Sport Today|||0|0|General Sports|News and results from around the world.
BBC News|1463965200|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463967000|The Week in Parliament|20/05/2016||0|0|General News,Current Affairs|A round-up of the week's proceedings in Parliament, presented by Alicia McCarthy.
BBC News|1463968800|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463970600|Dateline London|21/05/2016||0|0|reserved|Foreign correspondents currently posted to London look at events in the UK through outsiders' eyes, and at how the issues of the week are being tackled around the world.
BBC News|1463972400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463974200|HARDtalk|23/05/2016||0|0|Interview|Interviews with newsmakers and personalities from across the globe.
BBC News|1463976000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463977800|World Business Report|22/05/2016||0|0|General Social,Political Issues,Economics|The latest business news, with informed analysis.
BBC News|1463978700|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1463979600|Breakfast|||0|0|General Social,Political Issues,Economics|Round-up of national and international news, plus the latest from the money markets.
BBC News|1463988600|BBC Business Live|23/05/2016||0|0|General News,Current Affairs|A look at the global business stories.
BBC News|1463990400|Victoria Derbyshire|23/05/2016||0|0|News Magazine,Current Affairs|Daily news and current-affairs programme offering discussion of breaking stories, exclusive interviews and audience interaction via social media.
BBC News|1463997600|BBC Newsroom Live|23/05/2016||0|0|General News,Current Affairs|A chance to stay up to date on the day's leading stories, with the latest breaking news as it happens.
BBC News|1464004800|BBC News at One; Weather|23/05/2016||0|0|News|
BBC News|1464006600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464008400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464012000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464015600|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464019200|BBC News at Five|23/05/2016||0|0|News|The BBC News at Five O'Clock with in-depth discussions and analysis as well as breaking news.
BBC News|1464022800|BBC News at Six; Weather|23/05/2016||0|0|News|
BBC News|1464024600|Sportsday|||0|0|General Sports|Results and analysis from countrywide events.
BBC News|1464025500|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464026400|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464030000|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464031800|HARDtalk|23/05/2016||0|0|Interview|Interviews with newsmakers and personalities from across the globe.
BBC News|1464033600|Outside Source|||0|0|reserved|
BBC News|1464035400|Outside Source|||0|0|reserved|
BBC News|1464037200|BBC News at Ten|23/05/2016||0|0|News|
BBC News|1464039000|Sportsday|||0|0|General Sports|Results and analysis from countrywide events.
BBC News|1464039900|The Papers|23/05/2016 - 1||0|0|reserved|No need to wait until tomorrow morning to see what's in the papers - tune in to BBC News and hear a lively, informed and engaging conversation about the next day's papers.
BBC News|1464040800|BBC News|||0|0|News|The latest national and international stories as they break.
BBC News|1464041700|Sportsday|||0|0|General Sports|Results and analysis from countrywide events.
BBC News|1464042600|The Papers|23/05/2016 - 2||0|0|reserved|No need to wait until tomorrow morning to see what's in the papers - tune in to BBC News and hear a lively, informed and engaging conversation about the next day's papers.
BBC News|1464043500|Meet The Author|||0|0|reserved|Writers talk about their latest books.
BBC News|1464044400|Newsday|||0|0|News Magazine,Current Affairs|
BBC News|1464046200|HARDtalk|23/05/2016||0|0|Interview|Interviews with newsmakers and personalities from across the globe.(n)
BBC News|1464048000|Newsday|||0|0|News Magazine,Current Affairs|
BBC News|1464049800|Asia Business Report|23/05/2016||0|0|News Magazine,Current Affairs|Live from Singapore the essential business news as it breaks and a look ahead to the news that will shape the business day.(n)
BBC News|1464050700|Sport Today|||0|0|General Sports|News and results from around the world.(n)
BBC News|1464051600|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464053400|Monday in Parliament|23/05/2016||0|0|General News,Current Affairs|Highlights of the day's proceedings in Parliament.(n)
BBC News|1464055200|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464057000|Reporters|21/05/2016||0|0|reserved|A weekly showcase of the best reports from the BBC's global network of correspondents.(n)
BBC News|1464060600|HARDtalk|24/05/2016||0|0|Interview|Interviews with newsmakers and personalities from across the globe.(n)
BBC News|1464062400|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464064200|World Business Report|23/05/2016||0|0|General Social,Political Issues,Economics|The latest business news, with informed analysis.(n)
BBC News|1464065100|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464066000|Breakfast|||0|0|General Social,Political Issues,Economics|Round-up of national and international news, plus the latest from the money markets.(n)
BBC News|1464075000|BBC Business Live|24/05/2016||0|0|General News,Current Affairs|A look at the global business stories.(n)
BBC News|1464076800|Victoria Derbyshire|24/05/2016||0|0|News Magazine,Current Affairs|Daily news and current-affairs programme offering discussion of breaking stories, exclusive interviews and audience interaction via social media.(n)
BBC News|1464084000|BBC Newsroom Live|24/05/2016||0|0|General News,Current Affairs|A chance to stay up to date on the day's leading stories, with the latest breaking news as it happens.(n)
BBC News|1464091200|BBC News at One; Weather|24/05/2016||0|0|News|
BBC News|1464093000|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464094800|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464098400|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464102000|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464105600|BBC News at Five|24/05/2016||0|0|News|The BBC News at Five O'Clock with in-depth discussions and analysis as well as breaking news.(n)
BBC News|1464109200|BBC News at Six; Weather|24/05/2016||0|0|News|
BBC News|1464111000|Sportsday|||0|0|General Sports|Results and analysis from countrywide events.(n)
BBC News|1464111900|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464112800|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464116400|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464118200|HARDtalk|24/05/2016||0|0|Interview|Interviews with newsmakers and personalities from across the globe.(n)
BBC News|1464120000|Outside Source|||0|0|reserved|
BBC News|1464121800|Outside Source|||0|0|reserved|
BBC News|1464123600|BBC News at Ten|24/05/2016||0|0|News|
BBC News|1464125400|Sportsday|||0|0|General Sports|Results and analysis from countrywide events.(n)
BBC News|1464126300|The Papers|24/05/2016||0|0|reserved|No need to wait until tomorrow morning to see what's in the papers - tune in to BBC News and hear a lively, informed and engaging conversation about the next day's papers.(n)
BBC News|1464127200|BBC News|||0|0|News|The latest national and international stories as they break.(n)
BBC News|1464128100|Newsnight|24/05/2016||0|0|News Magazine,Current Affairs|Analysis of the day's events, presented by Emily Maitlis.(n)
BBC Parliament|1463893200|Select Committees|||0|0|General Social,Political Issues,Economics|Recorded coverage of the work of committees set up to investigate aspects of public policy and society.
BBC Parliament|1463913000|The Week in Parliament|20/05/2016||0|0|General News,Current Affairs|A round-up of the week's proceedings in Parliament, presented by Alicia McCarthy.
BBC Parliament|1463914800|America This Week|||0|0|General Education,Science|Highlights of the week in politics in the USA from C-SPAN.
BBC Parliament|1463918400|Washington Journal|||0|0|General Social,Political Issues,Economics|Highlights of the week from the USA.
BBC Parliament|1463925600|The Wales Report|The Wales Report with Huw Edwards||0|0|General Social,Political Issues,Economics|With five weeks until the referendum on Britain's membership of the EU, the broadcaster examines what impact an in or out vote will have on farming in Wales. Plus, the latest from the Senedd with Felicity Evans.
BBC Parliament|1463927700|The View|||0|0|General Social,Political Issues,Economics|Mark Carruthers presents a review of the week's political news, including reports on the latest events at Stormont and Westminster. Plus, comment and analysis with studio guests.
BBC Parliament|1463930100|Sunday Politics Scotland|22/05/2016||0|0|General Social,Political Issues,Economics|The week's events at Westminster, presented by Andrew Neil, with Andrew Kerr reporting from around Scotland. Also includes the day's news headlines.
BBC Parliament|1463932500|Sunday Politics Northern Ireland|22/05/2016||0|0|General Social,Political Issues,Economics|The week's events at Westminster with Andrew Neil and reports from around the Province with Mark Carruthers, plus the day's news headlines.
BBC Parliament|1463934000|Sunday Politics Wales|22/05/2016||0|0|General Social,Political Issues,Economics|The week's events at Westminster presented by Andrew Neil and reports from around Wales with Arwyn Jones, plus the day's news headlines.
BBC Parliament|1463935500|BOOKtalk|||0|0|General Arts,Culture|Mark D'Arcy presents a discussion of publications relating to the world of politics, including interviews with authors and commentators.
BBC Parliament|1463936400|Question Time|||0|0|Discussion,Debate|David Dimbleby chairs the debate from Walsall in the West Midlands, where the panel comprises Conservative Energy Secretary Amber Rudd, Labour former Cabinet Minister Yvette Cooper, Liberal Democrat leader Tim Farron, Ukip deputy leader Paul Nuttall and broadcaster Paul Mason.
BBC Parliament|1463940000|The Andrew Marr Show|22/05/2016||0|0|General News,Current Affairs|The political journalist presents a round-up of the week's stories, interviewing key figures and leafing through the Sunday papers.
BBC Parliament|1463943600|Select Committees|||0|0|General Social,Political Issues,Economics|Recorded coverage of the work of committees set up to investigate aspects of public policy and society.
BBC Parliament|1463958000|Sunday Politics London|22/05/2016||0|0|News Magazine,Current Affairs|The week's events at Westminster, presented by Andrew Neil. Including news and a regional round-up.
BBC Parliament|1463962500|Political Highlights|||0|0|General Social,Political Issues,Economics|Recorded coverage of political and parliamentary highlights.
BBC Parliament|1463979600|Westminster Hall|||0|0|General Education,Science|Recorded coverage of House of Commons proceedings in Westminster Hall from Thursday 19 May.
BBC Parliament|1463990400|The Week in Parliament|20/05/2016||0|0|General News,Current Affairs|A round-up of the week's proceedings in Parliament, presented by Alicia McCarthy.
BBC Parliament|1463992200|Select Committees|||0|0|General Social,Political Issues,Economics|Recorded coverage of the work of committees set up to investigate aspects of public policy and society.
BBC Parliament|1464010200|House of Commons|Live House of Commons: 23/05/2016||0|0|General Education,Science|Live coverage of the day's proceedings in the House of Commons.
BBC Parliament|1464040800|Monday in Parliament|23/05/2016||0|0|General News,Current Affairs|Highlights of the day's proceedings in Parliament, presented by Joanna Shinn.
BBC Parliament|1464042600|Lords Questions|23/05/2016||0|0|General Social,Political Issues,Economics|Recorded coverage of questions in the House of Lords.
BBC Parliament|1464044400|Daily Politics|23/05/2016||0|0|Discussion,Debate|Parliamentary proceedings interspersed with discussions, interviews and reports from correspondents around the country. Presented by Jo Coburn.(n)
BBC Parliament|1464048000|House of Lords|||0|0|General Social,Political Issues,Economics|Recorded coverage of Monday's business in the House of Lords.(n)
BBC Parliament|1464076800|Monday in Parliament|23/05/2016||0|0|General News,Current Affairs|Highlights of the day's proceedings in Parliament, presented by Joanna Shinn.(n)
BBC Parliament|1464078600|Select Committees|Live Select Committees||0|0|General Social,Political Issues,Economics|Live coverage of the work of committees set up to investigate aspects of public policy and society.(n)
BBC Parliament|1464085800|House of Commons|Live House of Commons: 24/05/2016||0|0|General Education,Science|Live coverage of the day's proceedings in the House of Commons.(n)
BBC Parliament|1464114600|House of Lords|Live House of Lords: 24/05/2016||0|0|General Social,Political Issues,Economics|Live coverage of the day's proceedings in the Palace of Westminster.(n)
BBC Parliament|1464127200|Tuesday in Parliament|24/05/2016||0|0|General News,Current Affairs|Highlights of the day's proceedings in Parliament, presented by Alicia McCarthy.(n)
BBC Parliament|1464129000|Lords Questions|24/05/2016||0|0|General Social,Political Issues,Economics|Recorded coverage of questions in the House of Lords.(n)
Channel 4|1463879100|Hollyoaks|||0|0|Soap,Melodrama|Omnibus. Scott is infuriated that he has been duped by Mercedes, while Pete is furious when Cleo tries to delay their plans, leaving her conflicted between her heart and her head. Elsewhere, Silas and Lindsey break into the Roscoes' house.
Channel 4|1463886600|The Three Day Nanny|||2|1|Documentary|Professional nanny Kathryn Mewes restores order to more households in distress, starting with the Morrisen family in Newbury. Mum Laura and three-year-old son Frankie are constantly at odds with each other, and the youngster's behaviour is tearing his parents apart. After moving in, Kathryn implements her own three-day action plan to help them sort out their problems.
Channel 4|1463889900|Posh Pawnbrokers|||1|8|Antiques,Collectibles|At Nikolas Patrick pawnbrokers in Kent, brothers Charlie and Patrick receive an Olympic torch that the owner wants £10,000 for, as well as some designer bags and a collection of antique firearms. Love is in the air for a newly engaged couple in Sheffield, and some rare footwear comes in.
Channel 4|1463892900|Salvage SOS|||1|1|Documentary|Documentary following an American architectural salvage crew, who recover historically important features from buildings due to be demolished so they can be incorporated into restoration projects. Salvagers Robert Kulp and Mike Whiteside visit Izard Farmhouse in Copper Hill, Virginia, and remove a bay window, a stairwell, a stove and vintage poplar wood, and deliver a Victorian doorway to its new home.
Channel 4|1463894400|Salvage SOS|||1|3|Documentary|The crew goes looking for salvage in the Robert E Lee Hotel, a six-storey establishment in Lexington, Virginia, that was built in 1926. The team emerges with a sink, subway-style tiles, a pair of French doors and some 1920s urinals. Plus, making a coffee table from a salvaged panel and some old printing plates and a search for vintage finds in a junkyard.
Channel 4|1463895900|Salvage SOS|||1|4|Documentary|The team goes looking for salvage in a grist mill in Virginia that was built in 1905, coming out with patina doors, granite mill stones and running gears. Plus, the guys also make a bar out of Egyptian iron and wood and buy a 1950s exercise machine.
Channel 4|1463897400|The King of Queens|Female Problems||2|2|Sitcom|Carrie becomes close friends with the new neighbour, leaving a jealous Doug feeling unwanted. American comedy set in New York, starring Kevin James.
Channel 4|1463898900|The King of Queens|Assaulted Nuts||2|3|Sitcom|Doug tries to get out of going to the bank with Carrie, claiming he is too busy at work, but a stapler-inflicted injury in a delicate area makes him see the error of his ways. Comedy, starring Kevin James.
Channel 4|1463900400|Frasier|Visions of Daphne||6|22|Sitcom|Daphne agrees to marry Donny, but has a vision that suggests he is wrong for her, and tempts fate by turning to Niles for advice on how to proceed.
Channel 4|1463902200|Frasier|Shut Out in Seattle - Part One||6|23|Sitcom|Part one of two. Daphne's engagement to Donny leaves Niles feeling down, so he seeks solace in the arms of a younger woman. Frasier keeps getting his girlfriend's name wrong, Martin's relationship with Bonnie turns sour, and Roz cannot bring herself to break up with Bulldog.
Channel 4|1463904000|Frasier|Shut Out in Seattle - Part Two||6|24|Sitcom|Part two of two. Niles and Roz take extreme action to solve dilemmas in their respective love lives. Comedy, starring Kelsey Grammer, David Hyde Pierce and Peri Gilpin.
Channel 4|1463905800|Sunday Brunch|||5|14|Cooking|Tim Lovejoy and Simon Rimmer are joined by guests wildlife presenter Steve Backshall, comedian James Acaster and actress Maddy Hill.
Channel 4|1463916600|Step Up||2006|0|0|General Movie,Drama|An aspiring ballerina finds her life turned upside down when she encounters a troubled street-smart teenager from the wrong side of town. But as the pair get together to work on a dance project, they develop a mutual admiration, and love begins to blossom between them. Romantic drama, starring Channing Tatum and Jenna Dewan. Edited for language and violence.
Channel 4|1463923800|Evolution||2001|0|0|Adventure|Two science teachers investigate a mysterious meteor and discover it is oozing a strange fluid containing millions of minuscule but rapidly evolving organisms - which start to turn into terrifying alien monsters with a taste for human flesh. Sci-fi comedy, starring David Duchovny, Orlando Jones, Julianne Moore, Seann William Scott, Dan Aykroyd and Ted Levine. Edited for language.
Channel 4|1463931000|Location, Location, Location|Lake District and Scottish Highlands Revisits||23|1|Property|House-hunting show with Kirstie Allsopp and Phil Spencer. The property experts catch up with two couples who hoped to realise dreams of finding a new home and business. Catherine and Mark wanted to move from the Midlands to the Lake District with plans to set up a hot-tub company, while Christine and Keith gave up life in Cambridgeshire to go in search of a hotel to run in the Highlands.
Channel 4|1463934600|A Place in the Sun: Winter Sun|||0|0|Tourism,Travel|Jasmine Harman helps a couple find a new home in the Mar Menor area of the the Costa Calida, where they hope to have a sea view and space to hold barbecues.
Channel 4|1463938200|Channel 4 News|22/05/2016||0|0|General Sports|Including sport and weather.
Channel 4|1463940000|Penelope Keith's Favourite Villages|||0|0|Documentary|The actress travels around Britain visiting villages in different parts of the country, and discovers how people's attitudes have changed to these small communities. Her trip takes her to villages in Devon, Cornwall, Scotland and the Lake District, with the help of insights from the illustrated 1930s Batsford Guides.
Channel 4|1463943600|The Best Exotic Marigold Hotel||2011|0|0|Comedy|Seven English pensioners looking for a fresh start are drawn to an advert for a hotel in the Indian city of Jaipur, and plan to spend their retirement there. They arrive to find the building dilapidated but are won over by the enthusiastic young manager, and each embarks on their own adventures in the city. Comedy drama, starring Judi Dench, Bill Nighy, Maggie Smith and Dev Patel. Edited for language.
Channel 4|1463952300|Gogglebox|||7|14|General Show,Game Show|The nation's favourite armchair critics share their opinions on what they have been watching during the week. The programme captures their instant reactions and lively - sometimes emotional - discussions from the comfort of their own homes.
Channel 4|1463956200|Hitchcock||2012|0|0|Biopic|Fact-based drama about the making of Alfred Hitchcock's Psycho. The film-maker is forced to fund the controversial project personally in the face of disinterest from the studios, while the financial strain and his lecherous behaviour begin to take their toll on his relationship with wife and creative partner Alma Reville. Starring Anthony Hopkins, Helen Mirren and Scarlett Johansson.
Channel 4|1463962500|Come Dine with Me|Hertfordshire||11|46|Challenge,Reality Show|Amir Hezarah kicks off the dinner parties in Hertfordshire, with a strategy to be on his best behaviour for the first night, before turning into his `real self' for the rest of the week. He is confident of impressing his guests with an Iranian feast of lamb stew and rose-water ice-cream.
Channel 4|1463964300|Come Dine with Me|Hertfordshire||11|47|Challenge,Reality Show|Cleanliness fanatic Claire Diamond hosts the second dinner party in Hertfordshire, hoping to impress with a menu of crispy chilli chicken, roast rack of lamb with potato dauphinoise and a large dessert of pana cotta, meringue and chocolate cheesecake. However, as the evening unfolds the simplicity of the menu upsets one of the guests and a shocking discovery is made in the bathroom.
Channel 4|1463966100|Come Dine with Me|Hertfordshire||11|48|Challenge,Reality Show|Would-be pop star Charles Maximilian Winnington Leftwich hosts the third dinner party in Hertfordshire, featuring an elaborate menu and an outdoor music performance. Unfortunately, it is not an easy ride for him as his guests struggle with his starter and rain threatens to spoil the barbecue.
Channel 4|1463967600|Come Dine with Me|Hertfordshire||11|49|Challenge,Reality Show|Diane Mitham hosts the penultimate dinner party in Hertfordshire. She hopes to impress with a menu of carrot and coriander soup, chicken lemon drizzle and witches' deadly cream scoop, and the evening gets off to an interesting start when she introduces her beloved pet - an eight-year-old tarantula.
Channel 4|1463969400|Come Dine with Me|Hertfordshire||11|50|Challenge,Reality Show|Hairdresser Mel Steel hosts the final day of the competition in Hertfordshire, and demonstrates her culinary skills with a mix of French and Caribbean dishes. The guests are shocked by her request for them to arrive in fancy dress, leaving her hopes of winning the £1,000 prize resting on the merits of her eclectic menu.
Channel 4|1463971200|Win It Cook It|||1|21|General Show,Game Show|Simon Rimmer and guest judge Matt Tebbutt compare chicken and meatball dishes.
Channel 4|1463972700|Location, Location, Location|Liverpool||17|4|Property|Kirstie Allsopp and Phil Spencer head to Liverpool, where they help two women with their house-hunting. Veronica Wright is a mother of two teenage boys, while Catherine Callaghan plans to set up a therapy business at home, so the experts face a tough challenge bringing the women's different lifestyles together under one roof. Student Kate Harland also receives advice on how to get on the property ladder.
Channel 4|1463976300|Fifteen to One|||0|0|Game Show,Quiz|Sandi Toksvig hosts the general knowledge quiz, in which 15 contestants are pitted against one another in the hope of securing a place in the end-of-series final when a £40,000 jackpot will be up for grabs.
Channel 4|1463979600|Countdown|20/05/2016||0|0|Game Show,Quiz|Nick Hewer and Rachel Riley present the words-and-numbers game, with journalist and broadcaster Janet Street-Porter in Dictionary Corner.
Channel 4|1463982300|Will & Grace|Something Borrowed, Someone's Due||4|18|Sitcom|Part two of two. The duo struggle to adjust to life in their new apartment and resort to devious means to get their old home back - but everything is put on hold when Ellen goes into labour. Comedy, starring Eric McCormack, Debra Messing and Leigh-Allyn Baker.
Channel 4|1463983800|Will & Grace|Cheatin' Trouble Blues||4|19|Sitcom|Will is so glad to hear his parents have settled their differences that he treats them to a cruise for their forthcoming anniversary, but is shocked to discover the pair have secrets to hide. Blythe Danner and Sydney Pollack guest star.
Channel 4|1463985300|Everybody Loves Raymond|Tasteless Frank||9|12|Sitcom|Frank puts salt on Marie's home-made lasagne, causing her to think she is turning into a terrible cook, but Ray and Robert discover their father has lost his sense of taste - apparently because of a potency medication he is taking. Comedy, starring Peter Boyle, Doris Roberts, Ray Romano and Brad Garrett.
Channel 4|1463986800|Everybody Loves Raymond|Sister-in-Law||9|13|Sitcom|Amy chats non-stop through a basketball game, and Ray responds by suggesting to Robert that she talks too much - a criticism she does not take well. Comedy, starring Monica Horan and Ray Romano.
Channel 4|1463988600|Everybody Loves Raymond|The Power of No||9|14|Sitcom|Debra cannot understand why Ray keeps turning down her advances - not realising that playing it cool is all part of his latest devious plan to get what he wants. Comedy, starring Ray Romano.
Channel 4|1463990400|Frasier|Momma Mia||7|1|Sitcom|Martin and Niles meet the new woman in Frasier's life - and discover to their surprise that she looks just like his mother. Comedy, guest starring Rita Wilson (Sleepless in Seattle), alongside Kelsey Grammer, John Mahoney and David Hyde Pierce.
Channel 4|1463992200|Frasier|Father of the Bride||7|2|Sitcom|Martin and Frasier inadvertently offer to pay for Daphne's wedding, while Niles sinks into gloom as the marriage approaches and tries to console himself by dating someone new - unaware she is a prostitute. Comedy, starring Kelsey Grammer.
Channel 4|1463994000|Frasier|Radio Wars||7|3|Sitcom|The station shock-jocks decide to play practical jokes - and Frasier's pompous manner makes him the ideal target for their dubious humour. Starring Kelsey Grammer and David Hyde Pierce.
Channel 4|1463995800|Undercover Boss Canada|||3|4|Documentary|General manager Gail Souter and operations manager Kristine Hubbard go undercover in their own privately owned taxi company - Beck Taxi. The mother-and-daughter team mingles with the workforce to learn more about the problems its drivers face.
Channel 4|1463999400|Four in a Bed|||7|16|General Show,Game Show|The contest begins at the Black Lion in Halland, East Sussex, where host Nigel Fright gets off to a shaky start when a kettle goes missing from one of the rooms. Later, he takes the guests to a salsa class, where Sherrill Tacy and Hayley Cotton are surprised by some of his dance moves.
Channel 4|1464001200|Channel 4 News Summary|24/05/2016||0|0|News|Includes news headlines and weather.
Channel 4|1464001500|Four in a Bed|||7|17|General Show,Game Show|The competition moves to the Wheatsheaf Inn in Exning, near Newmarket, Suffolk, where guests are welcomed by owner Ken Clutterbuck and employee Ginny Trow. The proprietor tries to win his rivals round with his unique sense of humour, but tensions rise when the contestants go for a spin on a go-kart track.
Channel 4|1464003300|Four in a Bed|||7|18|General Show,Game Show|Sherrill Tacy hosts at the Sherwood Guest House in New Brighton on the Wirral, and is praised for the establishment's value for money. However, there is upset when her breakfast leaves a lot to be desired, and her final review is far from perfect.
Channel 4|1464005100|Four in a Bed|||7|19|General Show,Game Show|Final hosts Mark and Rachael Dann welcome the contestants to the Big Bear Lodge in Shropshire. They face the tough job of trying to keep the rift between some of the guests to a minimum in their ski-themed B&B, and their afternoon activity of canoeing raises a few laughs but accusations of cheating occur when the boys begin to get competitive.
Channel 4|1464007200|Four in a Bed|||7|20|General Show,Game Show|The contestants featured throughout the week reunite to revisit the highs and lows of their various stays, and as the B&B owners confront their critics face to face, they discover what the rival parties really thought of the quality of service that they encountered. After the deliberations are over, the winning guest house is announced.
Channel 4|1464009000|Fifteen to One|||5|24|Game Show,Quiz|Sandi Toksvig hosts the general knowledge quiz, in which 15 contestants are pitted against one another in the hope of securing a place in the end-of-series final when a £40,000 jackpot will be up for grabs.
Channel 4|1464012600|Countdown|||0|0|Game Show,Quiz|Nick Hewer and Rachel Riley host the long-running words-and-numbers game, with Michael Buerk joining Susie Dent in Dictionary Corner.
Channel 4|1464015600|Couples Come Dine with Me|||2|43|Cooking|The doubles-version of the culinary challenge series heads to North Devon, where busy parents Matt and Sarah are the first hosts, but their decision to serve crisps as canapes does not go down well with some of their rivals. Next up are competitive `foodies' James and Laura, who put together a similar menu to their predecessors - but with more flair. The final party is thrown by am-dram couple Jake and Ian, and their guests' have high expectations that the pair's mushroom bruschetta starter and casserole main look set to miss.
Channel 4|1464019200|Four in a Bed|||14|36|General Show,Game Show|The competition begins at the Cuban-inspired Brovey Lair in Ovington, Norfolk, where owners Mike and Tina Pemberton kick things off with a salsa class, much to the horror of Sam Millidge and Nathan Pearce. Next morning, the open-plan restaurant and breakfast room causes issues for Richard and Sheryl Middleton, while Tina and Mike aren't happy with their feedback.
Channel 4|1464021000|Shipping Wars UK|||2|16|Documentary|Shahbaz transports a giant rat sculpture made of scrap metal and junk to the set of an indie movie in Bedford, while Laurie takes two converted shipping container homes from Newquay, Cornwall, to Manchester.
Channel 4|1464022800|The Simpsons|The Bob Next Door||21|22|Animated Movie,Drama|A new neighbour moves in next door to the family and proves popular with everyone - but Bart is convinced he is actually Sideshow Bob in disguise and sets out to unmask his arch-enemy. With the guest voice of Kelsey Grammer.
Channel 4|1464024600|Hollyoaks|||0|0|Soap,Melodrama|Scott organises a fairy light surprise for John Paul at The Folly, but he is overcome by guilt about Sally. Sienna feels under pressure, and elsewhere, Darren places bets on how long Trevor and Grace's marriage will last.
Channel 4|1464026400|Channel 4 News|24/05/2016||0|0|General Sports|Including sport and weather.
Channel 4|1464029700|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Vote Leave campaign.
Channel 4|1464030000|Eating Well with Hemsley + Hemsley|||1|3|Cooking|Even though Jasmine and Melissa Hemsley eat a diet totally free from gluten and grain, they still love baking and this edition features a selection of recipes for healthy living. After stocking up on alternatives to flour such as ground almonds and coconut flour, they make cinnamon banana bread that is perfect for breakfast, and gingernut cookies ideal for an afternoon snack. Always on the lookout for substitutes for refined sugar, the sisters visit two urban beekeepers in London who make raw honey.
Channel 4|1464031800|Food Unwrapped|||8|3|General Education,Science|Jimmy Doherty heads to the Spanish city of Seville to look for the mysterious ingredient that gives marmalade its bitter tang, while Kate Quilton meets an entrepreneur who has developed an ecosystem that could revolutionise the future of fish farming. Matt Tebbutt hits the streets to see how billy goat meat goes down with the British public.
Channel 4|1464033600|24 Hours in A&E|||11|2|Medicine,Health|Train driver Andy, 48, is rushed in after falling 12ft from a tree while cutting branches and landing on his feet, badly fracturing both ankles, and doctors are concerned the impact may have caused life-changing damage to critical nerves and blood vessels in his feet and legs. Angela, 59, has come to St George's as her heart has been beating at over 150bpm for eight hours, risking stroke and other complications. Cardiologist Dr Arun's attempts to bring down her pulse using a powerful drug aren't successful, so he decides to electrically shock her heart to reset it.
Channel 4|1464037200|Very British Problems|||2|3|Comedy|Famous faces offer their views on issues faced while on holiday, talking about those bizarre behaviours Brits display when they're out of our comfort zone and bombarded with languages, customs and situations they just don't understand Grace Dent and Alex Brooker share their airport taxi abduction anxieties, while other topics raised include how to stop holiday friendships with other Brits developing and the collective sigh of relief when it's all over. With contributions by James Corden, Jack Whitehall, David Tennant, Catherine Tate, Danny Dyer, Vic Reeves and Bob Mortimer. Last in the series.
Channel 4|1464041100|8 Out of 10 Cats Does Countdown|||7|9|Comedy|Jimmy Carr hosts the words-and-numbers panel game, with Sean Lock and guest captain Joe Wilkinson joined by Seann Walsh and Danny Dyer. Susie Dent is in Dictionary Corner, receiving a helping hand from Bill Bailey, while Rachel Riley looks after the numbers and letters.
Channel 4|1464044700|Random Acts|||0|0|General Arts,Culture|Eric Wareheim showcases more creative short films, including animations by the This Is It Collective and artists Kyle Platts and Andy Baker. An evocative snapshot of life in Huddersfield is set to music in Lucy Luscombe's video for electronic music duo Darkstar and there's an art film shot in the Balkans by Gery Georgieva for Friez.(n)
Channel 4|1464046500|24 Hours in Police Custody|The Black Balaclava||4|5|Documentary|The Bedfordshire police look into a rash of armed robberies in Luton, all of which have one thing in common - the victims were threatened at knifepoint. With no decent CCTV images to positively identify the two suspects who remain at large, the police need to fall back on some good old-fashioned detective skills.(n)
Channel 4|1464050100|Ramsay's Kitchen Nightmares USA|Hot Potato Cafe||3|1|Cooking|The chef again comes to the aid of failing American restaurants, starting in Fishtown, Philadelphia, where he tries to help the three owners of the Hot Potato Cafe, which has not made a profit in two years. Spurred on by a scathing review by an influential critic, he makes radical changes to alter the staff's attitudes and create food that is up to his own exacting standards.(n)
Channel 4|1464053100|The World's Most Extreme|Runways||1|5|General Education,Science|An exploration of the most unusual airports on the planet, including a runway squeezed between skyscrapers, a landing strip carved into mountains and an airport where the runway disappears with every tide. Plus, a military base that has been under repeated attacks for 10 years.(n)
Channel 4|1464056400|Posh Pawnbrokers|||1|7|Antiques,Collectibles|In Sheffield, London Road Pawnbrokers boss Dan hunts for a local artist regarding potentially valuable paintings, and an unusual silver sombrero could be worth a small fortune.(n)
Channel 4|1464059700|Kirstie's Fill Your House for Free|||0|0|DIY|Kirstie Allsopp stocks a Glasgow shop with furniture that has been sourced for free, transforming the items then offering them to people to furnish their homes.(n)
Channel 4|1464060900|Win It Cook It|||1|22|General Show,Game Show|The cooks compete for ingredients including crab meat and ricotta, and try to avoid fish heads and lime pickle, by answering the most questions correctly, before creating dishes for the enjoyment of host Simon Rimmer and guest chef Tony Singh.(n)
Channel 4|1464062700|Location, Location, Location|South-East London||17|1|Property|Two pairs of buyers enlist the help of Kirstie Allsopp and Phil Spencer to find their ideal properties in south-east London. Cruise ship workers Peter and Jason are looking forward to setting up home together in the popular suburb of Beckenham, while designers Nadine and Toby want a house in need of refurbishment within their £350,000 budget.(n)
Channel 4|1464066000|Countdown|||0|0|Game Show,Quiz|Nick Hewer and Rachel Riley host the long-running words-and-numbers game, with Michael Buerk joining Susie Dent in Dictionary Corner.(n)
Channel 4|1464068700|Will & Grace|Went to a Garden Potty||4|20|Sitcom|Will brings home the last remaining memento of his parents' marriage - an ugly garden gnome that he and his brothers bought them for their anniversary. Meanwhile, Jack worries about being typecast in heterosexual roles. Eric McCormack and Sean Hayes star.(n)
Channel 4|1464070200|Will & Grace|He Shoots, They Snore||4|21|Sitcom|Will accompanies Elliot to a basketball tournament after Jack drops out at the last minute, while Grace has a hard time teaching a design class to students with a short attention span. Eric McCormack and Debra Messing star.(n)
Channel 4|1464071700|Everybody Loves Raymond|Pat's Secret||9|15|Sitcom|Pat asks Robert to keep her cigarette habit a secret - but he later has to come up with an excuse when Amy smells smoke on him, leading to a string of revelations for the family.(n)
Channel 4|1464073200|Everybody Loves Raymond|Finale||9|16|Sitcom|In the last-ever episode of the American comedy, Ray has a brush with death while undergoing minor surgery, but pulls through - leaving his family uncertain over whether to tell him what happened.(n)
Channel 4|1464075000|Everybody Loves Raymond|Pilot||1|1|Sitcom|A chance to see the pilot episode of the comedy series. Debra tires of having to deal with Ray's interfering mother, grumpy father and resentful brother, who constantly show up out of the blue, and a white lie has embarrassing consequences. Starring Ray Romano and Patricia Heaton.(n)
Channel 4|1464076800|Frasier|Everyone's a Critic||7|4|Sitcom|Niles takes a new position as a magazine art critic, prompting a jealous Frasier to respond by launching his own arts show. Comedy, starring Kelsey Grammer and David Hyde Pierce.(n)
Channel 4|1464078600|Frasier|The Dog That Rocks the Cradle||7|5|Sitcom|Martin returns from a friend's funeral upset by how it was conducted, and begins to plan his own memorial. Meanwhile, sacked DJ Bulldog takes the opportunity to embark on an entirely new career - in pizza delivery. Comedy, starring Kelsey Grammer.(n)
Channel 4|1464080400|Frasier|Rivals||7|6|Sitcom|Niles and Frasier fall out, each convinced the other is secretly coveting his date. Comedy, starring Kelsey Grammer and David Hyde Pierce.(n)
Channel 4|1464082200|Undercover Boss Canada|||4|2|Documentary|Richard Andersen, the new CEO of sports and entertainment complex Northlands, is seeking to turn around the company's fortunes - so he goes undercover to find out what his employees make of his changes. He dons a fat suit and a new identity, and soon makes discoveries about staff morale and equipment, before the story of one worker's loss makes him realise the important steps he has to take.(n)
Channel 4|1464085800|Four in a Bed|||7|21|General Show,Game Show|The contest begins at One4 B&B in Cheltenham, where debonair art-dealing host Nick Purchase hopes to prove his that his establishment offers the best value for money. However, things get off to a less-than-ideal start when a life-drawing class leaves one of his guests in a fit of nervous giggles.(n)
Channel 4|1464087600|Channel 4 News Summary|24/05/2016||0|0|News|Includes news headlines and weather.(n)
Channel 4|1464087900|Four in a Bed|||7|22|General Show,Game Show|The competition moves to the Windy Bottom B&B in Maidstone, Kent, where owners Gloria Barnett and Dave Goulding try to impress their guests with a trip to Leeds Castle. However, a proprietor manages to offend one of her rivals, and another is not impressed at being allocated a Versace-themed room.(n)
Channel 4|1464089700|Four in a Bed|||7|23|General Show,Game Show|The third visit is to the Jolly Carter pub in Bolton, Greater Manchester, run by Phil and Angie Sutcliffe. Despite a few nerves about the accommodation not measuring up, the room inspections go well, but the guests' verdict on the afternoon's roller disco remains to be seen.(n)
Channel 4|1464091500|Four in a Bed|||7|24|General Show,Game Show|John Humberstone hosts at the 18-room Alexandra Hotel in Llandudno, where he hopes the scaffolding on the outside of his establishment will not ruin his chances. However, when one of the guests gets locked in a bathroom and there is a slip-up with towels and teabags, it seems he has plenty of other things to worry about.(n)
Channel 4|1464093600|Four in a Bed|||7|25|General Show,Game Show|The contestants featured on the show reunite to revisit the highs and lows of their various stays, and as the B&B owners confront their critics face to face, they discover what the rival parties really thought of the quality of service that they encountered. After the deliberations are over, the winning guest house is announced.(n)
Channel 4|1464095400|Fifteen to One|||5|25|Game Show,Quiz|Sandi Toksvig hosts the general knowledge quiz, in which 15 contestants are pitted against one another in the hope of securing a place in the end-of-series final when a £40,000 jackpot will be up for grabs.(n)
Channel 4|1464099000|Countdown|24/05/2016||0|0|Game Show,Quiz|Nick Hewer and Rachel Riley host as contestants race against the clock to pit their wits against vowels, consonants and numbers. Michael Buerk is in Dictionary Corner with Susie Dent.(n)
Channel 4|1464102000|Couples Come Dine with Me|||2|1|Cooking|Three couples from Leeds compete to host the best dinner party, beginning with construction manager Martin and his wife Amanda, who are determined to win. They are rivalled by competitive engaged couple Amy and Nico who impress with their entertainment and Hannah and Nick, who try to prove their doubters wrong by cooking duck to order.(n)
Channel 4|1464105600|Four in a Bed|||14|37|General Show,Game Show|The competition moves on to its second Norfolk B&B of the week, The Orangery, where Ricky and Vicky Kerrison's guests get competitive at an outdoor activity centre and try to leap from as high as possible on a jumping tower. Perfectionist Richard loses his nerve while young Sam and Nathan race to the top, and Vicky is determined to take them on.(n)
Channel 4|1464107400|Shipping Wars UK|||2|17|Documentary|Dave and Jenny head to Shrewsbury to deliver a giant aquarium that weighs 700kg. The 87 mile trip from Leicester involves a detour via Solihull to pick up some aggressive tropical fish.(n)
Channel 4|1464109200|The Simpsons|The Ten-Per-Cent Solution||23|8|Animated Movie,Drama|Things look bleak for Krusty the Clown when his TV show is binned and he is dropped by his talent agency. But then he is reunited with the veteran agent (Joan Rivers) who got him started in showbusiness all those years ago, and together they plan his big comeback.(n)
Channel 4|1464111000|Hollyoaks|||0|0|Soap,Melodrama|Grace is furious that her tyres have been slashed and tells Darren to replace them, only to find his betting book and the bets he has been taking on her wedding. Meanwhile, James talks John Paul into spending the day with him.(n)
Channel 4|1464112800|Channel 4 News|24/05/2016||0|0|General Sports|Including sport and weather.(n)
Channel 4|1464116100|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|A referendum broadcast by the Stronger in Europe campaign, ahead of the Referendum on the United Kingdom's membership of the European Union, on June 23rd.(n)
Channel 4|1464116400|Obsessive Compulsive Cleaners|Obsessive Compulsive Country House Cleaners||7|2|Documentary|Cleaners Kelly from County Durham and Dave from Surrey move into Forcett Hall in North Yorkshire. Owners James and Alison want to open a B&B, but with the bedrooms piled to the rafters with junk and vines growing through the windows, they and son Will are going to need all the help they can get transforming the Georgian manor into a des res once more.(n)
Channel 4|1464120000|How to Get a Council House|||4|3|Documentary|Cameras follows those who have come to the UK from abroad and have no option but to turn to the council for housing. They include Florin, his wife and their five children who have relocated from Romania for a better life in Britain but, without a home or a job, they face the prospect of having to sleep rough. Viewers also meet Monika from Poland and her Ugandan husband Frederick who have fallen behind on their rent and are now facing eviction.(n)
Channel 4|1464123600|Britain's Weirdest Council Houses|||0|0|Documentary|Tenants who have gone the extra mile to turn their local authority lodgings into unique homes, and the surprising stories behind each transformation. They include the painter-decorator who turned his Brighton terrace into a replica of the Sistine Chapel, and the pensioner who spent decades recreating the interior of a merchant navy ship in his flat on the 11th floor of a Portsmouth tower block.(n)
Channel 4|1464127500|24 Hours in A&E|||11|2|Medicine,Health|Train driver Andy, 48, is rushed in after falling 12ft from a tree while cutting branches and landing on his feet, badly fracturing both ankles, and doctors are concerned the impact may have caused life-changing damage to critical nerves and blood vessels in his feet and legs. Angela, 59, has come to St George's as her heart has been beating at over 150bpm for eight hours, risking stroke and other complications. Cardiologist Dr Arun's attempts to bring down her pulse using a powerful drug aren't successful, so he decides to electrically shock her heart to reset it.(n)
More4|1463872800|8 Out of 10 Cats Does Countdown|||4|4|Comedy|Jimmy Carr hosts the comedy panel show's version of the words-and-numbers game, with team captains Sean Lock and Jon Richardson joined by guests Jason Manford and Stephen Mangan. Tim Key joins Susie Dent in Dictionary Corner, while Joe Wilkinson causes trouble for Rachel Riley at the board.
More4|1463876700|Father Ted|Speed 3||3|3|Sitcom|Dougal takes over as Craggy Island's new milkman, but his predecessor, local womaniser Pat Mustard, returns to exact an explosive revenge on Ted for getting him sacked. Starring Ardal O'Hanlon and Dermot Morgan.
More4|1463878800|Father Ted|The Mainland||3|4|Sitcom|Dougal and Ted visit the mainland, where they bump into actor Richard Wilson - and discover the hard way that he does not take kindly to being confused with his comic alter ego Victor Meldrew. Dermot Morgan and Ardal O'Hanlon star.
More4|1463880600|Blue Eyes|The Wake||1|9|Adult Movie,Drama|Trapped with Mattias at the Veritas hideout, Sofia tends to his wounds, but an unsettling feeling torments her: Elin is contacted by an unexpected party who suggests a collaboration that could benefit them both, while the police identify Gustav through the CCTV pictures from the stock exchange. Thriller, starring Karin Franz Korlof and Adam Lundgren. In Swedish.
More4|1463903700|River Cottage Bites|||0|0|Cooking|Short highlights from Hugh Fearnley-Whittingstall's adventures at the smallholding, revealing the secrets to whipping up simple culinary treats.
More4|1463905500|Jamie's 15 Minute Meals|Fish Stew and Asian Beef||1|2|Cooking|Jamie Oliver continues to present quick and easy recipes. In this edition, he prepares flashy fish stew with saffron sauce and garlic bread, before making seared Asian beef, best noodle salad and ginger dressing.
More4|1463907300|A Place in the Sun: Home or Away|Nottingham v Barcelona||5|9|Property|Jason and Inge are torn over whether to buy a new home in Nottingham or start afresh in Barcelona, so appeal to Jonnie Irwin and Jasmine Harman for advice. The experts find affordable properties in both places, hoping the house-hunters will finally be able to make up their minds.
More4|1463911200|Homes by the Med|||1|5|General Arts,Culture|Charlie Luxton heads to the Costa del Sol, where he meets a couple who have built an extraordinary modern home that is designed like a cruise ship, but on dry land.
More4|1463914800|Come Dine with Me|Manchester||3|56|Challenge,Reality Show|Interior designer Carlos Buller kicks off a series of dinner parties in Manchester and impresses his guests with his unusual flat. However, a dispute with budding artist Karen Oulton threatens his chance of winning the £1,000 prize at the end of the week.
More4|1463916900|Come Dine with Me|Manchester||3|57|Challenge,Reality Show|Susan Brickell, a housing officer who has never thrown a formal dinner party before, hosts the second dinner party in Manchester. She aims to serve holiday-inspired Greek fare, but nerves get the better of her. To make matters worse, she is suffering from a hangover following the previous night's get-together.
More4|1463918700|Come Dine with Me|Manchester||3|58|Challenge,Reality Show|Performance artist and vegetarian Dan Cumberland prepares three curries and a dal in the hope of winning the £1,000 prize when he hosts the third night of the competition in Manchester. Stuart Burke throws his saffron tea away while the host is not looking, but is surprisingly won over by the main course. However, problems arise when it comes to serving the kulfi dessert, which is frozen solid.
More4|1463920800|Come Dine with Me|Manchester||3|59|Challenge,Reality Show|Contemporary artist Karen Oulton tries to claw her way back into her fellow contestants' good books by conjuring up an international feast for her dinner party in Manchester. However, she quickly manages to upset nightclub manager Stuart Burke with her strategy of preparing a four-course meal, when everyone else is cooking three.
More4|1463922600|Come Dine with Me|Manchester||3|60|Challenge,Reality Show|Nightclub manager Stuart Burke hosts the final meal of the week in Manchester, and hopes to secure the top prize with an inspired modern British menu. The evening gets off to a promising start as the food lover serves cocktails to his guests, but takes a turn for the worse when an argument ends in tantrums and tears.
More4|1463924400|Four in a Bed|||13|16|General Show,Game Show|The contest begins at Pauline Cox's Wharfe House in Wetherby, West Yorkshire, and a visit to a local vineyard sees a clash between guest Mike Hepker and Tash Thorne.
More4|1463926500|Four in a Bed|||13|17|General Show,Game Show|The B&B owners visit Wortwell Hall Barn in Norfolk, run by husband-and-wife duo Clive and Jenny Aylett, but when the pair's rivals arrive, Pauline Cox and Claire Smith have difficulty locating their favourite appliance. Publicans Mike Pearce and Tash Thorne are astonished to discover they cannot lock their room's door. In the morning, some of the guest make awkward requests to change their breakfast orders, causing professional chef Clive to experience a meltdown in the kitchen that leads to a fundamental error.
More4|1463928600|Four in a Bed|||13|18|General Show,Game Show|The contestants travel to Bath Lodge Castle in Somerset for the third day of the competition, where they are wowed by Karen and Mike Hepker's luxury castle experience. Although the guests are disappointed at the bathroom fixtures and fittings, they are given the chance to vent their emotions during an afternoon of painting in the castle grounds. Plus, tensions rise between Mike and Tash at dinner, and harsh comments at feedback lead the hosts to suspect game playing.
More4|1463930400|Four in a Bed|||13|19|General Show,Game Show|The final visit of the week is to The Old Lodge Hotel in Gosport, Hampshire, run by publicans Mike Pearce and Tash Thorne. Karen Hepker is disappointed with the honeymoon suite, while Clive and Jenny Aylett find a dubious looking splash guard in the shower. A boat tour backfires when Jenny struggles with her water phobia and at dinner Karen takes the opportunity to tell the others exactly what she thinks of them. But things really kick off when it comes to feedback time.
More4|1463932200|Four in a Bed|||13|20|General Show,Game Show|Wharfe House hosts Pauline Cox and Claire Smith begin a bitter debate, demanding to know why their beds caused such a sleepless night. Accusations subsequently fly in all directions and walk-outs look on the cards as tensions mount leading to the payments being revealed.
More4|1463934300|Come Dine with Me|York||19|31|Challenge,Reality Show|Training guru Steve Carlyle hosts the first party in York, but a sophisticated evening, complete with a butler, does nothing to boost his reputation as he competes to win the £1,000 prize at the end of the week.
More4|1463936100|Come Dine with Me|York||19|32|Challenge,Reality Show|Trevor Rooney, who leads tours of supposedly haunted sites in York, hosts the second dinner party in the city at a bric-a-brac warehouse. He also has several spooky surprises in store for his guests, including a magic show, a paranormal-themed menu and a ventriloquist's doll that spends the evening flirting with the female diners.
More4|1463937900|Come Dine with Me|York||19|33|Challenge,Reality Show|The third dinner party in York is hosted by Annie Albericci, who hopes to bring peace, love and harmony to the table with her festival-chic-themed evening. However, things go from bad to worse for Annie when the male guests find a racy photo of her.
More4|1463939700|Come Dine with Me|York||19|34|Challenge,Reality Show|Nurse Yvonne McGill hosts the fourth dinner challenge in York and goes for a 1960s-themed party, including a game of Snog, Marry, Avoid? and a Beatles tribute band. Meanwhile, guest Steve reveals his celebrity crush.
More4|1463941800|Come Dine with Me|York||19|35|Challenge,Reality Show|Foodie Rebecca Ryan hosts the final dinner party in York, and hopes to impress her guests by throwing a Hollywood-themed evening of glitz and glamour, before the winner of the £1,000 prize is announced.
More4|1463943600|Grand Designs New Zealand|||1|6|Property|Chris Moller meets a pastor and his wife who want a house with a perfect sea view, so take the step of building a three storey home on a crumbling cliff with a sheer drop below.
More4|1463947200|Ghost||1990|0|0|Fantasy|The spirit of a murdered executive tries to find a way to help his girlfriend bring his killer to justice and enlists the aid of a fraudulent medium - who is amazed and baffled when her psychic powers turn out to be all too real. Romantic fantasy, starring Patrick Swayze, Demi Moore, Tony Goldwyn and an Oscar-winning Whoopi Goldberg.
More4|1463956500|24 Hours in A&E|||2|14|Medicine,Health|A busy night shift sees a series of men admitted with various problems. Father-of-six Stacey is experiencing breathing difficulties, but his demanding attitude appears to mask a vulnerability. Twenty-year-old Sam is brought in after being attacked outside a nightclub and has possible injuries to the neck and spine. He is nervous because his father died at the hospital and, with a broken nose, is worried he may have lost his looks. Henry has an electrician's exam the following morning but has been hiccuping for three days. Registrar Faheem is determined to diagnose the problem and get him well in time.
More4|1463960100|24 Hours in A&E|||3|1|Medicine,Health|Documentary following life inside one of Britain's busiest A&E departments at King's College Hospital in south London. A doctor is shocked when a young woman arrives in resus with life-threatening swelling on her brain following a random attack by a stranger on the streets, while a mother faces an agonising wait as tests are carried out on her 12-year-old son, who was hit by a car and airlifted to King's by emergency medics. A 90-year-old former circus performer is also in A&E after collapsing at home, and news of his colourful past quickly circulates among the staff.
More4|1463964000|Father Ted|The Passion of St Tibulus||1|3|Sitcom|Bishop Brennan orders Ted and Dougal to campaign against a controversial film - but as a result of their protest it becomes the biggest box-office hit in Craggy Island's history. Comedy, starring Dermot Morgan, Ardal O'Hanlon, Frank Kelly and Pauline McLynn.
More4|1463966100|Father Ted|Competition Time||1|4|Sitcom|TV personality Henry Sellers arrives to judge an all-priest version of Stars in Their Eyes, prompting intense rivalry between the star-struck Craggy Island clerics and their Rugged Island counterparts. Comedy, with Dermot Morgan.
More4|1463968200|Grand Designs New Zealand|||1|6|Property|Chris Moller meets a pastor and his wife who want a house with a perfect sea view, so take the step of building a three storey home on a crumbling cliff with a sheer drop below.
More4|1463990100|Jamie's 15 Minute Meals|Chicken Fajitas and King Prawns||1|26|Cooking|Jamie Oliver prepares a selection of dishes including sizzling chicken fajitas, grilled peppers, salsa, rice and beans, plus prawn cocktail, king prawns and sun-dried pan bread.
More4|1463992500|A Place in the Sun: Winter Sun|Gran Canaria||4|0|Tourism,Travel|Jasmine Harman helps married couple Ali and Ben Brown from Kent find their ideal property abroad, as she shows them five places on the Spanish island of Gran Canaria.
More4|1463996400|The Long Gray Line||1955|0|0|Factual|A rebellious Irish immigrant to America does not initially fit in when he joins the army, but an instructor sees his potential as a teacher and takes him on as an assistant. He spends the next five decades at a military academy, becoming an inspirational figure to generations of soldiers through both World Wars. Fact-based drama, starring Tyrone Power and Maureen O'Hara.
More4|1464006300|Time Team|Lost Mines of Lakeland||20|6|Archaeology|Tony Robinson and the team head to the Lake District to look for copper, a forgotten piece of the nation's industrial heritage. There are nearly two dozen old mines across the mountains, some thought to have been established 400 years ago when the valleys would have been studded with workshops, scaffolding and water-powered machines, home to a brave band of Tudor miners. The team battles the rain, wind and dangerously unstable trackways, but the combination of sheer effort and hi-tech kit enables the experts to access the heart of an old mine.
More4|1464010200|Time Team|Horseshoe Hall||20|7|Archaeology|The team heads to the small county of Rutland to visit Oakham Castle, the most well-preserved 12th-century building in Britain. It was once home to the Norman knight Walkelin de Ferrers, who fought alongside Richard the Lionheart in the Crusades, and before that the residence of several Saxon kings and queens. Tony and the crew investigate de Ferrers' long-lost private quarters, but it takes three days of twists and turns to determine what the site looked like 900 years ago. To mark the visit, they also cast a giant Time Team horseshoe to add to the collection that has decorated the castle hall for half a millennium.
More4|1464014100|A Place in the Sun: Winter Sun|Gran Canaria||4|0|Tourism,Travel|Jasmine Harman helps married couple Ali and Ben Brown from Kent find their ideal property abroad, as she shows them five places on the Spanish island of Gran Canaria.
More4|1464018000|A Place in the Sun: Winter Sun|Mojacar||4|13|Tourism,Travel|London-based couple Rena Sodhi and Donna Carty want a second home they can escape to in Mojacar, southern Spain. Laura Hamilton finds a townhouse with stunning views for £25,000 less than their budget, but the buyers spot something even more tempting in the presenter's line up of possible purchases.
More4|1464021900|Selling Houses with Amanda Lamb|||2|5|Property|Homeowners in Leicester who are struggling to sell their properties receive help from the property expert to make their homes more appealing to buyer Panna, who has a budget of £275,000. Gurpal and Kiran need to inject some colour into their bland decor, while Sheetal could benefit from adding some furniture to her empty house, and Belinda and Spencer hesitate to make the recommended improvements.
More4|1464025800|George Clarke's Amazing Spaces|||4|2|General Education,Science|The architect meets a man trying to build the first UFO-styled prefabricated Futuro house seen in Britain for 50 years, and a woman creating a magical garden room using centuries-old techniques, involving earth, sand, straw and even human hair. George's Italian road trip takes him to a traditional old village, where he discovers the most modern of houses with an extraordinary design featuring a floating swimming pool. And, as he and Will get down to work on their wilderness retreat, there's a close shave involving an oak tree.
More4|1464029700|Grand Designs|||14|4|Property|Architect Patrick Bradley has come up with an unusual £100,000 house design built out of four 45ft shipping containers, welded together to form a giant cross and cantilevered over the top of a stream on the family farm in Co Derry. His mother is hoping the new home will help her son find a girlfriend, but the small budget and tight schedule soon pose problems. Kevin McCloud follows his progress.
More4|1464033600|The Supervet|||5|3|Vets,Pets|Professor Noel Fitzpatrick tends to a Newfoundland called Billy, who clocks up thousands of miles travelling back and forth from his home in Aberdeen for treatment on its legs. He also attempts to help Barney, a Yorkshire terrier that has a deformity in its neck that is compressing its spinal cord. For owners Linda and Barry, Noel is their last chance, but the operation involves high-risk surgery with no guarantee of success.
More4|1464037200|One Born Every Minute|||6|5|Family and Friends|Catherine and Simon went through years of fertility treatment to have their first son, which took a toll on their love life, but five years later, awaiting an elective C-section for their second baby, it's a different story - a spontaneous romantic evening resulted in an unexpected positive pregnancy test. Heather ran into complications during her first pregnancy and had to deliver twins at 24 weeks. They pulled through, but cerebral palsy and other issues have meant she is now a full-time carer to them both. She also has Alfie, and after he was born, she and partner Dan decided they would have a fourth child to give him a companion to help share the responsibility of siblings with a disability. Christian couple Naomi and Dan tied the knot young and had their first child 13 months ago. Now, they're back at Southmead for baby number two.
More4|1464041100|24 Hours in A&E|||3|2|Medicine,Health|Eighty-year-old Rose has fluid on her lungs and is having trouble breathing. Her daughters Christine, Sandra and Debbie put on brave faces around her bedside, convincing her that everything will be all right, but in the relatives' room there's high emotion as they contemplate life without their mother. Also in resus at King's College Hospital is Kevin, a 55-year-old trucker who has sustained injuries in a road accident.
More4|1464045000|Embarrassing Bodies|Thailand - Part One||5|1|General Education,Science|Dr Dawn Harper heads to Thailand with Dr James Logan, who infests himself with a parasitic hookworm as he investigates the ailments Britons could catch there. Back in the UK, Dr Pixie McKenna meets a woman with an addiction to coffee enemas, and Dr Christian Jessen advises a patient who has had breast enhancement surgery.(n)
More4|1464048900|The Supervet|||5|3|Vets,Pets|Professor Noel Fitzpatrick tends to a Newfoundland called Billy, who clocks up thousands of miles travelling back and forth from his home in Aberdeen for treatment on its legs. He also attempts to help Barney, a Yorkshire terrier that has a deformity in its neck that is compressing its spinal cord. For owners Linda and Barry, Noel is their last chance, but the operation involves high-risk surgery with no guarantee of success.(n)
More4|1464052800|One Born Every Minute|||6|5|Family and Friends|Catherine and Simon went through years of fertility treatment to have their first son, which took a toll on their love life, but five years later, awaiting an elective C-section for their second baby, it's a different story - a spontaneous romantic evening resulted in an unexpected positive pregnancy test. Heather ran into complications during her first pregnancy and had to deliver twins at 24 weeks. They pulled through, but cerebral palsy and other issues have meant she is now a full-time carer to them both. She also has Alfie, and after he was born, she and partner Dan decided they would have a fourth child to give him a companion to help share the responsibility of siblings with a disability. Christian couple Naomi and Dan tied the knot young and had their first child 13 months ago. Now, they're back at Southmead for baby number two.(n)
More4|1464056400|River Cottage Bites|||0|0|Cooking|River Cottage chef Gill Meller demonstrates how to make soft white rolls for lunchtime, and his colleague Gideon Hitchin presents a simple recipe for oatcakes.(n)
More4|1464076500|Jamie's 15 Minute Meals|Jerk Pork and Poached Chicken||1|10|Cooking|Chef Jamie Oliver prepares more quick meals, including his recipe for jerk pork with grilled corn and crunchy tortilla salad, as well as minestrone poached chicken and salsa verde.(n)
More4|1464078900|A Place in the Sun: Winter Sun|Mojacar||4|13|Tourism,Travel|London-based couple Rena Sodhi and Donna Carty want a second home they can escape to in Mojacar, southern Spain. Laura Hamilton finds a townhouse with stunning views for £25,000 less than their budget, but the buyers spot something even more tempting in the presenter's line up of possible purchases.(n)
More4|1464082800|Food Unwrapped|||2|1|General Education,Science|Jimmy Doherty, Matt Tebbutt and Kate Quilton travel the globe to explore the secrets behind mass-produced food. Jimmy visits cheese cellars in the south of France where mould is specially grown to be eaten, Kate is in Ukraine to discover which part of a chicken is used in a Kiev, while Matt finds out how shops sell English summer apples in the middle of winter.(n)
More4|1464084600|Hugh's 3 Good Things: Best Bites|||1|3|Cooking|Hugh Fearnley-Whittingstall creates a simple supper of clams, tomatoes and garlic.(n)
More4|1464085200|Please Sir||1971|0|0|Comedy|A put-upon teacher at an inner-city secondary school struggles to cope with his disruptive pupils and tempts fate by taking them on a fortnight's trip to an outdoor pursuits centre. Big-screen version of the TV comedy, starring John Alderton, Deryck Guyler, Noel Howlett, Joan Sanderson and Richard Davies.(n)
More4|1464092700|Time Team|Mystery of the Thames-side Villa||20|8|Archaeology|The experts head to a field in south Oxfordshire where significant findings were made by an inquisitive PhD student half a century ago, including a mosaic and the stone walls of a former Roman building. Tony Robinson and the crew examine aerial pictures showing clear building lines in the ground, and speak to the current landowner, a farmer who continues to uncover bricks and tiles. They try to evaluate the building's purpose and how the Thames may have shifted the remains over the course of two millennia.(n)
More4|1464096600|Time Team|The Lost Castle of Dundrum||20|9|Archaeology|Tony Robinson and the team search for the remains of a Norman castle in Dundrum, Co Down, one of Northern Ireland's most picturesque counties, exploring a territory established by renegade knight John de Courcy in the 12th century against the orders of King John. The castle was later rebuilt, and much of its replacement is still standing, but the experts are convinced that some of what remains dates from de Courcy's time - and discover that it may go back even further.(n)
More4|1464100500|A Place in the Sun: Winter Sun|Lanzarote||4|15|Tourism,Travel|Jasmine Harman helps couple Jane and David Turnbull, who have a budget of £80,000, to search for a house in Lanzarote. The property must have a lot of potential, and the pressure is on as it will eventually become their retirement home.(n)
More4|1464104400|A Place in the Sun: Winter Sun|Mar Menor||4|1|Tourism,Travel|Former pub landlady Janice Gibson wants to swap her Newcastle lifestyle for a new start in the Mar Menor area of southern Spain, so Laura Hamilton shows her a selection of properties starting from around £55,000.(n)
More4|1464108300|Selling Houses with Amanda Lamb|||2|6|Property|Three homeowners in Hucknall, Nottinghamshire, compete to sell their homes to first-time buyers George and Grace after making a number of improvements to their properties. Claire Michalski needs to complete some renovations, Claire Gadsby needs to de-clutter her abode, while Dave and his daughter Lauren add colour to their decor.(n)
More4|1464112200|George Clarke's Amazing Spaces|||4|3|General Education,Science|Will Hardie and George struggle to bring ancient Roman technology back to life and the build on their log cabin in the wilderness begins in earnest, while the road trip around Italy takes in an impressive fire station. The architect also meets David Moreton, a former Paralympic swimmer hoping to turn an old air ambulance into an amphibious crash pad for his charity fundraising tours, and DIY enthusiasts Ben and Michelle, who want to build a summerhouse for free, using hundreds of disused shipping pallets.(n)
More4|1464116100|Grand Designs|||14|6|Property|Natasha Cargill wants to build a home shaped like two enormous periscopes in rural Norfolk, but to obtain planning permission, she has to ensure not only that the materials are sustainable, but also agree to measure the transportation used to deliver them. If these strict criteria are not met, she won't be allowed to live there, and to add to the pressure, she has just £330,000 to spend on construction and six months to complete the project. Kevin McCloud follows her progress.(n)
More4|1464120000|Homes by the Med|||1|6|General Arts,Culture|Charlie Luxton travels to Puglia, Italy, and in the seaside town of Polignano a Mare, he visits a townhouse perched precariously over sea caverns. He also takes in a rural building in Alberbello with an unusual conical roof. Last in the series.(n)
More4|1464123600|999: What's Your Emergency|||2|3|Documentary|The documentary follows paramedics as they deal with mental-health cases. Maria Stanley is called to a multistorey car park, where she tries to talk a man away from the edge, while Kirsten Harper and Amy Siddall race to help a father who is having suicidal thoughts. In London, crews attend the scene of a failed suicide attempt that has left a middle-aged man trapped under a train.(n)
More4|1464127800|My Daughter the Teenage Nudist|||0|0|Documentary|Documentary following Mollie and Alex, who are part of a growing band of teenagers and twentysomethings who embrace the concept of public nudity away from designated places. Their aim is to normalise naturism and question the media's apparent obsession with perfect bodies. The programme asks why this lifestyle is gaining in popularity and finds out what parents think about their offspring revealing all in the most public of places.(n)
Film4|1463877600|Boomerang||1992|0|0|Comedy|A high-flying advertising executive is also an insatiable womaniser. However, he is brought down to earth with a bump by his glamorous new boss, who seduces him then breaks his heart, giving him a taste of the way he has previously treated women. Romantic comedy, starring Eddie Murphy, Robin Givens, Halle Berry, Grace Jones, Eartha Kitt and Chris Rock.
Film4|1463911200|Faintheart||2008|0|0|Comedy|Family man Richard finds solace from his humdrum life in the world of historical battle re-enactments. However, when his hobby sees him spend more time on the battlefield than at home, his wife leaves him for a gym instructor, forcing Richard to reassess his priorities. Romantic comedy, starring Eddie Marsan, Ewen Bremner, Jessica Hynes, Bronagh Gallagher, Tim Healy and Paul Nicholls.
Film4|1463918400|The Golden Compass||2007|0|0|Adventure|Orphan Lyra Belacqua lives in a parallel universe populated by magical and menacing characters. When her best friend becomes the latest in a long line of children to mysteriously vanish, she embarks on a perilous mission to uncover the dark secret behind their disappearance. Fantasy adventure based on Philip Pullman's novel Northern Lights, starring Dakota Blue Richards, Nicole Kidman, Daniel Craig and Eva Green. Featuring the voices of Ian McKellen, Kristin Scott Thomas and Kathy Bates.
Film4|1463926200|Marmaduke||2010|0|0|Comedy|An advertising executive tries to start a new life in California with his family and their lumbering, disaster-prone Great Dane. The friendly but clumsy dog accidentally causes chaos for his owners, until an incident at a surfing competition makes him a local celebrity. Comedy, with Lee Pace, and featuring the voice of Owen Wilson.
Film4|1463932500|Tooth Fairy||2010|0|0|Comedy|A minor-league ice hockey player is nicknamed the Tooth Fairy for knocking opponents' teeth out on the ice. When the cynical athlete discourages a young fan, he is forced to pay penance by spending a week as the real Tooth Fairy, rediscovering his dreams in the process. Family comedy, starring Dwayne Johnson, Ashley Judd, Stephen Merchant, Ryan Sheckler and Seth MacFarlane.
Film4|1463940000|Just Married||2003|0|0|Comedy|A newlywed couple are in for a rude awakening when they jet off on their dream honeymoon. They are looking forward to an enjoyable tour of Europe - but a series of chaotic events, plus the intervention of the bride's old flame, leaves them at each other's throats and their marriage in tatters. Romantic comedy, with Brittany Murphy, Ashton Kutcher, Christian Kane and David Moscow.
Film4|1463947200|The Hunger Games: Catching Fire||2013|0|0|Adventure|Katniss Everdeen's victory in a televised death match makes her a focus for revolution against the totalitarian nation she lives in. The rulers of the regime plot to crush dissent with a new series of games, in which past champions battle it out. Sci-fi adventure sequel based on the second book in Suzanne Collins' trilogy of novels, starring Jennifer Lawrence, Liam Hemsworth, Donald Sutherland and Philip Seymour Hoffman.
Film4|1463957400|House of Flying Daggers||2004|0|0|Adventure|Two imperial officers are sent to find the head of a rebel group, which threatens to destroy the Tang dynasty's tenuous grip on power. Their search leads the duo to a beautiful blind dancer, who they hope will take them to the mysterious and influential figure - but matters soon take an unexpected turn. Romantic period martial arts adventure from director Zhang Yimou, starring Zhang Ziyi, Takeshi Kaneshiro, Andy Lau and Song Dandan. In Mandarin.
Film4|1463965800|Kelly + Victor||2012|0|0|General Movie,Drama|Two strangers unhappy with their dull lives meet in a Liverpool nightclub and begin a purely sexual relationship that finally offers them the excitement they seek, while also providing them with an outlet for their darker urges. Drama based on Niall Griffiths' novel, starring Antonia Campbell-Hughes and Julian Morris.
Film4|1463997600|Hell in the Pacific||1968|0|0|War|An American GI and a Japanese soldier are marooned together on a deserted Pacific island during the Second World War. At first, the stranded pair are determined to kill each other, but as time passes they reach an impasse and realise they have to rely on each other to survive. Drama, starring Lee Marvin and Toshiro Mifune.
Film4|1464005100|Caprice||1967|0|0|Comedy|A cosmetics company employee goes undercover in a rival firm to try and steal the secret of their latest product - a miracle spray that keeps hair dry even underwater. Her assignment leads to a run-in with a secret agent, who is investigating something far more dangerous. Comedy thriller, starring Doris Day and Richard Harris.
Film4|1464012300|The Desert Fox||1951|0|0|War|German commander Rommel falls out of favour with Hitler following his defeat at El Alamein. On returning to his homeland, he is torn between his oath of loyalty and lack of faith in the Fuehrer's unstable leadership, prompting him to become involved in an assassination plot. Second World War drama, starring James Mason, Jessica Tandy, Cedric Hardwicke, Leo G Carroll and Luther Adler.
Film4|1464018600|The Man from Laramie||1955|0|0|Western|A cavalry officer determines to avenge the death of his brother, but rather than target the Apaches who killed him, he vows to go after the gang who supplied them with their weapons - leading to conflict with the sadistic son of an elderly rancher. Anthony Mann's Western, starring James Stewart, Arthur Kennedy, Donald Crisp and Cathy O'Donnell.
Film4|1464026100|Field of Dreams||1989|0|0|Fantasy|A farmer hears a mysterious voice inspiring him to mark out a baseball diamond in a cornfield - which, to his surprise, is visited by the ghost of the star player of the 1919 Chicago White Sox team, whose career was cut short by scandal. It later dawns on him the pitch has a greater purpose - to give people who have sacrificed important parts of their lives a second chance. Fantasy, starring Kevin Costner, Ray Liotta, Burt Lancaster and James Earl Jones.
Film4|1464033600|The Wolverine||2013|0|0|Adventure|The former member of the X-Men is lured out of hiding and travels to Japan, where a dying businessman offers him the chance to give up his immortality for a normal life. He ends up robbed of his superhuman powers by a mysterious scientist and is forced to protect the tycoon's granddaughter from a secret conspiracy's assassins. Superhero adventure spin-off, starring Hugh Jackman and Tao Okamoto.
Film4|1464042300|An Officer and a Gentleman||1982|0|0|General Movie,Drama|A Navy recruit undergoing officer training has an uneasy romance with a factory worker. He also attracts the attention of a tough, uncompromising sergeant, who sees his potential and is determined to push him to the limit. Romantic drama, starring Richard Gere, Debra Winger, Louis Gossett Jr, Robert Loggia, David Keith and David Caruso.
Film4|1464051300|Half Nelson||2006|0|0|General Movie,Drama|A teacher working in a tough inner-city school develops an addiction to crack cocaine. When a 13-year-old female student with a turbulent home life learns of his dependency, the discovery marks the beginning of an unlikely friendship between the pair. Drama, starring Ryan Gosling, Shareeka Epps and Anthony Mackie.(n)
Film4|1464084000|Footsteps in the Fog||1955|0|0|Historical,Period Drama|A prominent Victorian gentleman thinks he has got away with poisoning his wife, but his shrewd maid knows the sordid truth and uses it to blackmail him. As the killer's social standing improves, he realises he has to get rid of the scheming servant once and for all, but his plans to dispose of her lead him into even more danger. Period thriller, with Stewart Granger, Jean Simmons and Bill Travers.(n)
Film4|1464090300|Titanic||1953|0|0|Disaster Movie|An aristocratic woman flees her loveless marriage, taking her children with her and boarding the supposedly unsinkable ship as it embarks on its ill-fated maiden voyage. She is unaware her husband has followed her on board in an attempt to stop her leaving - but the pair's marital difficulties are soon overshadowed by the impending disaster. Drama, starring Clifton Webb, Barbara Stanwyck, Robert Wagner, Richard Basehart and Thelma Ritter.(n)
Film4|1464097500|Silent Running||1972|0|0|Science Fiction|A scientist, with the help of his three robot assistants, tends a huge garden aboard a space station, created to replenish an Earth ravaged by nuclear warfare. But his superiors' decision to abandon the project prompts him to embark on a desperate course of action. Ecological sci-fi drama, starring Bruce Dern, with Cliff Potts and Ron Rifkin.(n)
Film4|1464103800|The Lady Vanishes||1979|0|0|Mystery|An American heiress befriends an elderly lady on a continental train journey, but wakes one morning to find she has disappeared and the other passengers deny having ever seen the missing woman - leading to suspicions that a conspiracy is afoot. Remake of Hitchcock's 1938 mystery, starring Elliott Gould, Cybill Shepherd, Angela Lansbury, Herbert Lom, Arthur Lowe and Ian Carmichael.(n)
Film4|1464111000|Runaway Jury||2003|0|0|Literary Adaptation|A woman sets in motion a multimillion-dollar lawsuit against the manufacturer of the gun that was used to kill her husband - but her actions spark an unexpected series of events when a jury consultant for the defence tries to buy the verdict his clients want. Thriller, adapted from a novel by John Grisham, starring John Cusack, Gene Hackman, Dustin Hoffman, Rachel Weisz and Bruce Davison.(n)
Film4|1464120000|The Five-Year Engagement||2012|0|0|Comedy|A couple decide to get married, but before they can begin planning their wedding in earnest, a series of unforeseen events forces them to postpone the big day. As a career opportunity leads them to make a fresh start in another part of the country, second thoughts start to surface and the altar looks a very long way away. Romantic comedy, with Jason Segel, Emily Blunt and Rhys Ifans.(n)
Film4|1464128700|Predator 2||1990|0|0|Science Fiction|A Los Angeles cop, working to bring down the city's drug gangs, suspects Jamaican criminals when he discovers several of his targets killed and skinned alive. However, the culprit behind the murders reveals himself to be an alien big-game hunter - with the stealth and guile to outwit the police and criminals alike. Sci-fi sequel, starring Danny Glover, Bill Paxton, Gary Busey and Maria Conchita Alonso.(n)
ITV Anglia|1463872200|Jackpot247|||0|0|Game Show,Quiz|Viewers are offered the chance to participate in live interactive gaming from the comfort of their sofas, with an entertaining mix of roulette-wheel spins and lively chat from the presenting team. Featuring a variety of prizes and promotions.
ITV Anglia|1463882400|Murder, She Wrote|The Days Dwindle Down||3|21|Mystery|Jessica researches a 30-year-old murder case that may have led to the imprisonment of an innocent man. Starring Angela Lansbury and Richard Beymer.
ITV Anglia|1463885400|ITV Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV Anglia|1463893200|The Aquabats! Super Show|||0|0|Cartoons,Puppets|Action comedy following the fortunes of the Aquabats, a musical group of amateur superheroes.
ITV Anglia|1463894700|Pat & Stan|||0|0|Cartoons,Puppets|Animated fun with Pat the hippopotamus and Stan the dog.
ITV Anglia|1463895300|Dino Dan|||0|0|General Children's,Youth|Adventures for younger viewers following trainee paleontologist Dan Henderson and his friends.
ITV Anglia|1463895900|Dino Dan|||0|0|General Children's,Youth|Adventures for younger viewers following trainee paleontologist Dan Henderson and his friends.
ITV Anglia|1463896800|Signed Stories|Signed Stories: Share a Story||0|0|General Children's,Youth|A look behind the scenes of the Share a Story competition, meeting the competitors and the animators who turned their stories into short films.
ITV Anglia|1463897100|Sooty|||0|0|General Children's,Youth|Further adventures with ever-popular puppet pals Sooty, Sweep and Soo.
ITV Anglia|1463897700|Super 4|||0|0|Cartoons,Puppets|Animated comedy adventure series featuring a gang of heroes who protect the city of Technopolis and its King Kenric against evil elements.
ITV Anglia|1463898600|Nerds & Monsters|||0|0|Cartoons,Puppets|Animated comedy about a group of children exiled on an uncharted island, where they have to be smart if they are to survive relentless attacks by a tribe of hideous monsters.
ITV Anglia|1463899500|The Tom & Jerry Show|||0|0|General Children's,Youth|Madcap slapstick and mayhem as the celebrated cat and mouse plot against each other.
ITV Anglia|1463900400|Teen Titans Go|||0|0|Cartoons,Puppets|The teenage superheroes fight to save the world while getting up to mischievous antics.
ITV Anglia|1463901900|ITV News|||0|0|News|
ITV Anglia|1463902200|Weekend|||3|12|Talk Show|Aled Jones is joined by guests In the Club star Christine Bottomley and Supernanny's Jo Frost. Katherine Jenkins performs live in the studio and comedian Patrick Monahan provides his take on the latest news stories.
ITV Anglia|1463905500|Griff's Great Britain|Highlands||1|3|General Education,Science|Griff Rhys Jones explores the Highlands as he goes in search of Britain's second-largest bird of prey, travelling through the scenic and ancient landscape by a variety of means - but will he be able to track down the elusive golden eagle?.
ITV Anglia|1463907600|Peston on Sunday|||1|3|Discussion,Debate|Political magazine, presented by Robert Peston, with ITV News National Editor Allegra Stratton. Featuring reports on the latest issues and interviews with topical guests.
ITV Anglia|1463911200|FIA Formula E Championship|2016 Berlin ePrix Highlights||0|0|Motor Sport|The Berlin ePrix. Jennie Gow presents highlights of the eighth round of the season, staged on a track at the Alexanderplatz in the heart of the city. Lucas Di Grassi led the standings after seven rounds, with Britain's Sam Bird back in third place. With commentary by Jack Nicholls and Allan McNish, and reports from Nicki Shields.
ITV Anglia|1463914800|ITV News and Weather|||0|0|News|
ITV Anglia|1463915340|ITV Anglia Weather|||0|0|Weather|
ITV Anglia|1463915400|The Jeremy Kyle Show|22/05/2016 - 1||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.
ITV Anglia|1463919300|Planet's Got Talent|||1|4|Variety Show|Highlights from the Got Talent franchise around the world, featuring a man called Professor Splash who jumps into paddling pools from incredible heights, a Romanian who eats raw chicken, a parrot that speaks fluent English, a South Korean pensioner who picks a fight with a load of rocks, and a Chinese man performing one of the most dangerous acts ever seen on the show. Narrated by Warwick Davis.
ITV Anglia|1463921100|Fierce|Namibia||1|5|Wildlife|Naturalist Steve Backshall explores the wildlife in the landscapes of Namibia, southern Africa. He tracks two hungry cheetahs as they go on a hunt, stakes out a carcass to get up close to a group of vultures, and has a close encounter with an agitated lion as he helps a vet at work.
ITV Anglia|1463924700|Britain's Got Talent|||10|7|General Show,Game Show|Ant and Dec host the final round of auditions before the nationwide talent contest moves on to the next stage, the Judges' Decisions. One last selection of would-be stars demonstrate their signature skills to Simon Cowell, Alesha Dixon, Amanda Holden and David Walliams, in the hope of securing a place among the acts seeking a place in the semi-finals. However, there are no Golden Buzzers left to send promising stars straight through to the finals, so even the most eye-catching acts will have to fight for a place in the semi-finals.
ITV Anglia|1463929200|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1463930100|ITV News and Weather|||0|0|News|
ITV Anglia|1463931000|Live International Football|England v Turkey||0|0|Football - International|England v Turkey (Kick-off 5.15pm). Mark Pougatch presents coverage of the friendly encounter, which takes place at the Etihad Stadium in Manchester and serves as a Euro 2016 warm-up for both countries. This is the first time these sides have met since the qualifying campaign for Euro 2004, when two fiery games saw England claim a 2-0 home win and a 0-0 draw in Istanbul that secured their passage to Portugal. Roy Hodgson has already selected his squad for this summer's tournament in France, so he will be hoping the players can come through this encounter - and the upcoming friendlies with Australia and Portugal - with a clean bill of health. With analysis from Ian Wright and Lee Dixon, and commentary by Clive Tyldesley and Glenn Hoddle.
ITV Anglia|1463941800|Britain's Got Talent|Live Semi-Final||10|8|General Show,Game Show|Ant and Dec host the first semi-final of this year's contest. The audition process is complete, and has left judges Amanda Holden, David Walliams, Simon Cowell and Alesha Dixon with 45 acts to pick and choose from. Tonight, nine of them will be performing live in the hope of impressing both the panel and the TV audience. The winner of tonight's viewers' vote will automatically go through to the live grand final, before the two runners up face the judges to decide which of them will also win a place.
ITV Anglia|1463947200|Coronation Street|||0|0|Soap,Melodrama|Long-running drama with the residents of England's most famous cobbled street.
ITV Anglia|1463949000|Britain's Got Talent Results|Live Results||10|1|General Show,Game Show|Ant and Dec announce the results of tonight's viewers' vote to decide which act will make it through to the grand final. Judges Simon Cowell, David Walliams, Alesha Dixon and Amanda Holden will then select one of the runners up to join them. The show also features a performance by the cast of West End musical Motown.
ITV Anglia|1463950800|ITV News and Weather|||0|0|News|
ITV Anglia|1463951940|ITV Anglia Weather|||0|0|Weather|
ITV Anglia|1463952000|International Football Highlights|England v Turkey||0|0|Football - International|England v Turkey. Jacqui Oatley presents action from the friendly encounter, which took place at the Etihad Stadium in Manchester and served as a Euro 2016 warm-up for both countries. This was the first time these sides had met since the qualifying campaign for Euro 2004, when two fiery games saw England claim a 2-0 home win and a 0-0 draw in Istanbul that secured their passage to Portugal. Roy Hodgson has already selected his squad for this summer's tournament in France, so he will have been hoping the players would come through this encounter - and the upcoming friendlies with Australia and Portugal - with a clean bill of health. With analysis from Lee Dixon and Glenn Hoddle, and commentary by Clive Tyldesley.
ITV Anglia|1463955600|Premiership Rugby Union|2015/16 Semi-Finals||0|0|Rugby Union - Domestic|Mark Durden-Smith and David Flatman present highlights of the semi-finals, which were Saracens v Leicester Tigers at Allianz Park and Exeter Chiefs v Wasps at Sandy Park.
ITV Anglia|1463958900|Jackpot247|||0|0|Game Show,Quiz|Viewers are offered the chance to participate in live interactive gaming from the comfort of their sofas, with an entertaining mix of roulette-wheel spins and lively chat from the presenting team. Featuring a variety of prizes and promotions.
ITV Anglia|1463968800|Motorsport UK|2016 Donington Park||0|0|Motor Sport|Action from Donington Park, featuring the MSA Formula Championship and the Ginetta GT4 Supercup. Commentary by Richard John Neil.
ITV Anglia|1463971800|ITV Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV Anglia|1463976300|The Jeremy Kyle Show|22/05/2016 - 2||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.
ITV Anglia|1463979600|Good Morning Britain|23/05/2016||0|0|Magazine Show|A lively mix of news and current affairs, plus health, entertainment and lifestyle features.
ITV Anglia|1463988600|Lorraine|23/05/2016||0|0|General Education,Science|Entertainment and fashion news, as well as showbiz stories, cooking and celebrity gossip. Presented by Lorraine Kelly.
ITV Anglia|1463991900|The Jeremy Kyle Show|23/05/2016 - 1||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.
ITV Anglia|1463995800|This Morning|23/05/2016||0|0|General Education,Science|Phillip Schofield and Holly Willoughby present celebrity chat and lifestyle features, including a look at the stories making the newspaper headlines and a recipe in the kitchen. Including Local Weather.
ITV Anglia|1464003000|Loose Women|23/05/2016||0|0|Talk Show|Celebrity interviews and topical studio discussion from a female perspective.
ITV Anglia|1464006600|ITV Lunchtime News|||0|0|News|
ITV Anglia|1464008100|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1464008400|Judge Rinder|23/05/2016||0|0|General Education,Science|Cameras follow criminal barrister Robert Rinder as he takes on real-life cases in a studio courtroom.
ITV Anglia|1464012000|Dickinson's Real Deal|Prestatyn 2||12|0|General Show,Game Show|David Dickinson is in Prestatyn, north Wales, where experts Tony Geering, Corrie Jeffery and Stewart Hofgartner value items brought in by members of the public.
ITV Anglia|1464015540|ITV Anglia Weather|||0|0|Weather|
ITV Anglia|1464015600|Tipping Point|23/05/2016||0|0|Quiz Show|Game show, hosted by Ben Shephard, in which contestants answer questions to win turns on an arcade-style machine. Dropping tokens down a choice of four chutes, they hope to knock piles of them off a moving shelf - and the more they collect, the greater the prize fund. The player who has won the least amount is then eliminated, and the last one standing competes for a £10,000 jackpot.
ITV Anglia|1464019200|The Chase|||10|17|Quiz Show|Bradley Walsh presents as Steve, Virinder, Julie and Pat pit their wits against ruthless quiz genius the Chaser in the hope of winning a potential prize pot worth thousands of pounds. They work as a team and play strategically to answer general knowledge questions against the clock and race down the game board to the exit without being caught.
ITV Anglia|1464022800|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1464024300|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Vote Leave campaign.
ITV Anglia|1464024600|ITV Evening News|||0|0|News|
ITV Anglia|1464026400|Emmerdale|||0|0|Soap,Melodrama|Lawrence demands that Ronnie leave his family alone, only to find the plumber knows things he would rather keep secret. Doug tries to give Laurel a break from her worries, and Chrissie is delighted when her divorce comes through. Vanessa is less than thrilled when Carly invites Tracy to come and live with them, and Sam fears Megan is considering giving Jai another chance.
ITV Anglia|1464028200|Britain's Got Talent|Live Semi-final Two||10|9|General Show,Game Show|Ant and Dec present the second live semi-final, as nine more of the 45 chosen acts compete to impress judges Amanda Holden, David Walliams, Simon Cowell and Alesha Dixon and secure the all-important viewers' vote. At stake is the chance to appear at this year's Royal Variety Performance and win a life-changing cash prize of £250,000, with the act with the highest public vote going through automatically, while two runners-up fight it out for the judges' favour.
ITV Anglia|1464033600|Coronation Street|||0|0|Soap,Melodrama|With Johnny nowhere to be found, Roy offers to walk Carla down the aisle, but as she comes face to face with the groom, the bride tells Nick she wants to speak to him in private. Will the ceremony go ahead?.
ITV Anglia|1464035400|Britain's Got Talent Results|||10|2|General Show,Game Show|Ant and Dec announce the act with the highest number of public votes, automatically going through to the final. Simon Cowell, David Walliams, Amanda Holden and Alesha Dixon then decide which of the contestants in second and third place they want to see again. Plus, American pop-rock band One Republic perform.
ITV Anglia|1464037200|ITV News at Ten|23/05/2016||0|0|News|
ITV Anglia|1464039300|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1464039900|The Cube|Rhodri and Zoe||9|2|Game Show,Quiz|The high-pressure contest continues as Phillip Schofield invites more members of the public to step into the Cube for another selection of agility tests and skill trials that could see them score a jackpot of £250,000. This time, Welsh farmer Rhodri Jones hopes to win the cash prize to buy a prized bull, and barista Zoe Webster has her sights set on taking her family on a dream holiday.
ITV Anglia|1464043500|Murder, She Wrote|Time to Die||10|16|Mystery|Jessica is shocked to discover one of her writing students has been arrested on suspicion of murdering his stepfather, and makes a bid to help clear the boy's name. Angela Lansbury, Robert Beltran and Billy Gallo star.
ITV Anglia|1464046500|Jackpot247|||0|0|Game Show,Quiz|Viewers are offered the chance to participate in live interactive gaming from the comfort of their sofas, with an entertaining mix of roulette-wheel spins and lively chat from the presenting team. Featuring a variety of prizes and promotions.(n)
ITV Anglia|1464055200|The Jeremy Kyle Show|23/05/2016 - 2||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.(n)
ITV Anglia|1464058500|ITV Nightscreen|||0|0|General Education,Science|Text-based information service.(n)
ITV Anglia|1464062700|The Jeremy Kyle Show|23/05/2016 - 3||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.(n)
ITV Anglia|1464066000|Good Morning Britain|24/05/2016||0|0|Magazine Show|A lively mix of news and current affairs, plus health, entertainment and lifestyle features. Presented by Susanna Reid, Piers Morgan, Ben Shephard, Charlotte Hawkins and Sean Fletcher.(n)
ITV Anglia|1464075000|Lorraine|||0|0|General Education,Science|Director Jodie Foster talks about her latest film, Money Monster, which stars George Clooney and Julia Roberts. Presented by Lorraine Kelly.(n)
ITV Anglia|1464078300|The Jeremy Kyle Show|24/05/2016 - 1||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.(n)
ITV Anglia|1464082200|This Morning|24/05/2016||0|0|General Education,Science|Phillip Schofield and Holly Willoughby present celebrity chat and lifestyle features, including a look at the stories making the newspaper headlines and a recipe in the kitchen. Including Local Weather.(n)
ITV Anglia|1464089400|Loose Women|||19|0|Talk Show|Topical debate from a female perspective and celebrity interviews.(n)
ITV Anglia|1464093000|ITV Lunchtime News|||0|0|News|
ITV Anglia|1464094500|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1464094800|Judge Rinder|24/05/2016||0|0|General Education,Science|Cameras follow criminal barrister Robert Rinder as he takes on real-life cases in a studio courtroom.(n)
ITV Anglia|1464098400|Dickinson's Real Deal|Edinburgh 2||12|0|General Show,Game Show|David Dickinson and his team of dealers are in Edinburgh, where David Hakeney, Henry Nicholls and Helen Gardiner seek to pick more valuable items.(n)
ITV Anglia|1464101940|ITV Anglia Weather|||0|0|Weather|
ITV Anglia|1464102000|Tipping Point|24/05/2016||0|0|Quiz Show|Game show, hosted by Ben Shephard, in which contestants answer questions to win turns on an arcade-style machine. Dropping tokens down a choice of four chutes, they hope to knock piles of them off a moving shelf - and the more they collect, the greater the prize fund. The player who has won the least amount is then eliminated, and the last one standing competes for a £10,000 jackpot.(n)
ITV Anglia|1464105600|The Chase|||0|0|Quiz Show|Bradley Walsh presents as contestants Saroop, Karen, Milo and Natalie pit their wits against ruthless quiz genius the Chaser in the hope of winning a potential prize pot worth thousands of pounds. They work as a team and play strategically to answer general knowledge questions against the clock and race down the game board to the exit without being caught.(n)
ITV Anglia|1464109200|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1464110700|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Britain Stronger in Europe campaign.(n)
ITV Anglia|1464111000|ITV Evening News|||0|0|News|
ITV Anglia|1464112800|Emmerdale|||0|0|Soap,Melodrama|Lawrence is furious when Rakesh offers Ronnie a job overseeing the Mill conversion, and enlists Sam's help in a drastic attempt to get rid of him once and for all. Charity tries to frame Holly for stealing from Victoria's van, and a reluctant Jimmy is roped into keeping an eye on Ashley and Arthur - but ends up enjoying himself, and offers to help Doug with the secret supervision.(n)
ITV Anglia|1464114600|Britain's Got Talent|Live Semi-final Three||10|10|General Show,Game Show|Ant and Dec present the third live semi-final as more acts take to the stage in a bid to impress Simon Cowell, Alesha Dixon, David Walliams and Amanda Holden and reach the final. The victors will be in with a chance of scooping the £250,000 prize and a slot at the Royal Variety Performance.(n)
ITV Anglia|1464120000|Coronation Street|||0|0|Soap,Melodrama|With Jenny now guarding a captive Tracy for Johnny, it remains to be seen whether she will be able to escape and stop the wedding before it has even begun. How will Nick react to what Carla has to tell him?.(n)
ITV Anglia|1464121800|Britain's Got Talent Results|||10|3|General Show,Game Show|The viewers have spoken after another semi-final filled with talent, and the act with the highest number of votes goes straight through to the final. The two runners-up are then left at the mercy of the judges, who decide which of them deserves the remaining spot. Ant and Dec present, and guest Nick Jonas provides the music.(n)
ITV Anglia|1464123600|ITV News at Ten|24/05/2016||0|0|News|
ITV Anglia|1464125700|ITV News Anglia|||0|0|Regional News|
ITV Anglia|1464126300|Living with Quads|||0|0|Documentary|Any parent knows the challenges that a new baby brings, from the culture shock of nappy changes and sleepless nights to the realisation that time is no longer your own. Now imagine that multiplied by four. This one-off documentary follows the ups and downs of family life for people with quadruplets, meeting families with children of different ages - from babies to 10-year-olds - to reveal the joys, the occasional heartaches and the sacrifices that are necessary when a family expands by four overnight.(n)
ITV Anglia|1464129900|Columbo: A Stitch in Crime||1973|0|0|Police,Crime Drama|Surgeon Barry Mayfield decides he needs get rid of his colleague to speed along a research project. When his partner requires heart surgery, Mayfield performs the operation himself and discreetly arranges some fatal complications. However, when he also murders a nurse who suspects the truth, he attracts the attention of the slovenly sleuth. Crime drama, starring Peter Falk, Leonard Nimoy and Will Geer.(n)
ITV2|1463871900|Family Guy|Peter's Two Dads||5|10|Animated Movie,Drama|Peter discovers his mother had an affair while on holiday in Ireland 40 years previously, and crosses the Atlantic to search for his real father. Meanwhile, Stewie develops a love of punishment.
ITV2|1463873700|American Dad|Don't Look a Smith Horse in the Mouth||6|10|Animated Movie,Drama|Francine demands that Stan gives up his expensive SUV, so he buys a racehorse in a bid to win enough money to keep his petrol-guzzling car. Meanwhile, Steve enlists the aid of his friends to help an old acquaintance. Comedy, with the voices of Seth MacFarlane and Wendy Schaal.
ITV2|1463875500|American Dad|Shallow Vows||6|6|Animated Movie,Drama|Francine decides to drop her beauty regimen ahead of her 20th wedding anniversary, hoping to determine whether Stan loves her for more than her looks. However, the spy becomes upset that his wife has started to let herself go, and resorts to drastic measures when she asks him to renew their marital vows.
ITV2|1463877000|The Cleveland Show|Back to Cool||2|20|Animated Movie,Drama|Cleveland challenges Donna's ex-husband Robert to a Coolympics competition, hoping to prove his hip credentials to Cleveland Jr. Featuring the guest voice of Snoop Dogg.
ITV2|1463878500|The Cleveland Show|Your Show of Shows||2|21|Animated Movie,Drama|Rallo and his friends Bernard and Theodore perform in the school talent show, but their rap about fiscal responsibility proves unpopular with the student body. Meanwhile, Cleveland turns to daytime TV for answers when his own debut show is panned by critics. With the voices of Will.i.am and T-Pain.
ITV2|1463880000|@elevenish|||0|0|Comedy|Topical comedy series in which a cast of stand-ups, character actors and comedy groups share their thoughts on the past seven days through monologues, sketches and commentary.
ITV2|1463881200|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.
ITV2|1463892000|ITV2 Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV2|1463893200|Planet's Funniest Animals|||0|0|Nature,Animals|Humorous clips of pets and other animals in unusual situations.
ITV2|1463894400|Emmerdale|||0|0|Soap,Melodrama|Long-running soap following the ups and downs of village life amid the rolling scenery of the Yorkshire Dales.
ITV2|1463903700|Coronation Street|||0|0|Soap,Melodrama|Long-running drama with the residents of England's most famous cobbled street.
ITV2|1463913900|Take Me Out|||3|3|Game Show,Quiz|A personal trainer from Manchester, a football freestyler from Walsall, a Staffordshire student and a Bedford mobile-phone salesman enter the `love lift' in the hope of impressing 30 single women and winning a date - but must first get the female participants to keep their lights on as a sign of approval. Last week's couples go on their dates to discover whether they are a match made in heaven or hell. Paddy McGuinness presents.
ITV2|1463918400|A Little Princess||1995|0|0|Family|A wealthy English girl is sent to an austere New York boarding school, where she charms the other youngsters with her stories of life in India - until her father goes missing in action, leaving her destitute and in the hands of the wicked headmistress. Drama based on Frances Hodgson Burnett's classic novel, with Eleanor Bron, Liesel Matthews and Liam Cunningham.
ITV2|1463922300|FYI Daily|22/05/2016 - 1||0|0|News Magazine,Current Affairs|
ITV2|1463922600|A Little Princess||1995|0|0|Family|A wealthy English girl is sent to an austere New York boarding school, where she charms the other youngsters with her stories of life in India - until her father goes missing in action, leaving her destitute and in the hands of the wicked headmistress. Drama based on Frances Hodgson Burnett's classic novel, with Eleanor Bron, Liesel Matthews and Liam Cunningham.
ITV2|1463925300|The Smurfs 2||2013|0|0|Comedy|The tiny blue forest-dwelling creatures and their human friends go on a rescue mission to Paris. Their old foe Gargamel the evil wizard has created mischievous smurfs of his own and kidnapped Smurfette to learn the secret of her magic. Fantasy comedy sequel, starring Hank Azaria and Neil Patrick Harris, with the voices of Katy Perry and Christina Ricci.
ITV2|1463928900|FYI Daily|22/05/2016 - 2||0|0|News Magazine,Current Affairs|
ITV2|1463929200|The Smurfs 2||2013|0|0|Comedy|The tiny blue forest-dwelling creatures and their human friends go on a rescue mission to Paris. Their old foe Gargamel the evil wizard has created mischievous smurfs of his own and kidnapped Smurfette to learn the secret of her magic. Fantasy comedy sequel, starring Hank Azaria and Neil Patrick Harris, with the voices of Katy Perry and Christina Ricci.
ITV2|1463932500|Britain's Got Talent|||10|7|General Show,Game Show|Ant and Dec host the final round of auditions before the nationwide talent contest moves on to the next stage, the Judges' Decisions. One last selection of would-be stars demonstrate their signature skills to Simon Cowell, Alesha Dixon, Amanda Holden and David Walliams, in the hope of securing a place among the acts seeking a place in the semi-finals. However, there are no Golden Buzzers left to send promising stars straight through to the finals, so even the most eye-catching acts will have to fight for a place in the semi-finals.
ITV2|1463937300|Britain's Got More Talent|||10|7|General Show,Game Show|Stephen Mulhern hosts the companion show to the talent competition, going behind the scenes during the last round of auditions before the judges start to whittle down the successful candidates to their chosen semi-finalists.
ITV2|1463940900|Hulk||2003|0|0|Adventure|Scientist Dr Bruce Banner turns into the rampaging green Hulk after exposure to a huge dose of gamma radiation, prompting the military to embark on a no-holds-barred mission to destroy the monster. Meanwhile, Banner's unstable father resurfaces, holding the secret to his transformation. Comic-strip adventure from director Ang Lee, starring Eric Bana, Jennifer Connelly, Sam Elliott and Nick Nolte.
ITV2|1463944800|FYI Daily|22/05/2016 - 3||0|0|News Magazine,Current Affairs|
ITV2|1463945100|Hulk||2003|0|0|Adventure|Scientist Dr Bruce Banner turns into the rampaging green Hulk after exposure to a huge dose of gamma radiation, prompting the military to embark on a no-holds-barred mission to destroy the monster. Meanwhile, Banner's unstable father resurfaces, holding the secret to his transformation. Comic-strip adventure from director Ang Lee, starring Eric Bana, Jennifer Connelly, Sam Elliott and Nick Nolte.
ITV2|1463950800|Britain's Got More Talent|||10|8|General Show,Game Show|Stephen Mulhern goes behind the scenes of the talent competition's second live semi-final, featuring exclusive chats with celebrity guests, contestants and the judges.
ITV2|1463954400|Family Guy|Scammed Yankees||14|12|Animated Movie,Drama|Peter and Carter go to Africa to get their money back after they are swindled in an e-mail scam, while Brian pursues Meg's friend Patty.
ITV2|1463956200|Family Guy|It Takes a Village Idiot and I Married One||5|17|Animated Movie,Drama|Lois campaigns for election as mayor, but is only successful after dumbing down her political views to appeal to the electorate. However, the power of her office soon corrupts her and she begins to accept bribes to buy expensive things for herself. Meanwhile, Peter enjoys all the perks his status as `first lady' of Quahog brings him.
ITV2|1463958000|Family Guy|The Tan Aquatic with Steve Zissou||5|11|Animated Movie,Drama|An unfortunate experience on a tanning bed leaves Stewie convinced he has skin cancer. Meanwhile, Chris discovers rival paper boy Kyle has stolen one of his customers - so Peter beats him up.
ITV2|1463959800|American Dad|Brains, Brains and Automobiles||6|4|Animated Movie,Drama|Stan fears Francine will leave him if she realises how boring he is without Steve, Hayley and Roger in the house - so he concocts a scheme to have the alien move back in.
ITV2|1463961300|American Dad|Man in the Moonbounce||6|5|Animated Movie,Drama|Stan tries to live out the childhood he never had by playing pranks - but his adolescent adventures only succeed in landing him in jail - forcing Steve to become the man of the house.
ITV2|1463963100|The Cleveland Show|Hot Cocoa Bang Bang||2|22|Animated Movie,Drama|The family attends Comic-Con, where Cleveland plans to promote his creation Waderman. Meanwhile, Donna is horrified to discover that a blaxploitation film she starred in when she was younger is being screened at the event, and Cleveland Jr embarks on a mission to restore the annual gathering to its humble roots.
ITV2|1463964900|The Cleveland Show|BFFs||3|1|Animated Movie,Drama|Cleveland make an effort to bond with his friends by going on a camping trip, but the holiday takes a dangerous turn. Meanwhile, Donna encourages Rallo to prove he is as clever as his classmates by competing in a quiz tournament.
ITV2|1463966100|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.
ITV2|1463978700|ITV2 Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV2|1463979600|The Hot Desk|The Hot Desk: DNCE||0|0|General Music,Ballet,Dance|US band DNCE face a grilling over the Hot Desk.
ITV2|1463980200|Dinner Date|Jonathan||1|23|Cooking|Northampton bachelor Jonathan chooses three blind dates based on menus created by five potential partners. When the three dinners have been eaten, he decides who he wants to see again. Narrated by Charlotte Hudson.
ITV2|1463983200|The Ellen DeGeneres Show|||0|0|Talk Show|The host is joined by actor Alec Baldwin. Plus, a performance by Keith Urban with his song Wasted Time.
ITV2|1463986200|Emmerdale|||0|0|Soap,Melodrama|A social worker visits to see if Ashley is fit to look after Arthur, but he takes their agreement very badly. Lawrence asks Sam to sort out a leaking washing machine, but he unwittingly hires Ronnie Hale to do the job, forcing Chrissie to open up to Bernice. Jai refuses to take the hint that Megan is not interested in him, and Doug and Diane urge Pollard to throw Tracy out of the B&B.
ITV2|1463988000|Coronation Street|||0|0|Soap,Melodrama|Carla fears for her future with Nick after her plans to give him a stress-free day backfire, and Jenny flirts with Johnny at the factory and asks if he will give her a promotion. Meanwhile, Kevin arranges a summit in the hope that Izzy and Anna can settle their differences.
ITV2|1463989800|Coronation Street|||0|0|Soap,Melodrama|Nick is undecided about whether he can cope with moving to Devon and Izzy's revelation that she has been charged with possession of cannabis and assaulting a police officer causes amazement. Elsewhere, Jenny continues to play games with Johnny following her sewing lesson.
ITV2|1463991600|Psych|Dis-Lodged||2|14|Comedy|The duo investigate the death of a member of a local fraternity chaired by Lassiter's father-in-law. Comic detective drama, starring James Roday as a novice sleuth.
ITV2|1463994600|Britain's Got Talent|Live Semi-Final||10|8|General Show,Game Show|Ant and Dec host the first semi-final of this year's contest. The audition process is complete, and has left judges Amanda Holden, David Walliams, Simon Cowell and Alesha Dickson with 45 acts to pick and choose from. Tonight, nine of them will be performing live in the hope of impressing both the panel and the TV audience. The winner of tonight's viewers' vote will automatically go through to the live grand final, before the two runners up face the judges to decide which of them will also win a place.
ITV2|1464000300|Britain's Got Talent Results|Live Results||10|1|General Show,Game Show|Ant and Dec announce the results of tonight's viewers' vote to decide which act will make it through to the grand final. Judges Simon Cowell, David Walliams, Alesha Dixon and Amanda Holden will then select one of the runners up to join them. The show also features a performance by the cast of West End musical Motown.
ITV2|1464002100|Emmerdale|||0|0|Soap,Melodrama|A social worker visits to see if Ashley is fit to look after Arthur, but he takes their agreement very badly. Lawrence asks Sam to sort out a leaking washing machine, but he unwittingly hires Ronnie Hale to do the job, forcing Chrissie to open up to Bernice. Jai refuses to take the hint that Megan is not interested in him, and Doug and Diane urge Pollard to throw Tracy out of the B&B.
ITV2|1464003900|Coronation Street|||0|0|Soap,Melodrama|Carla fears for her future with Nick after her plans to give him a stress-free day backfire, and Jenny flirts with Johnny at the factory and asks if he will give her a promotion. Meanwhile, Kevin arranges a summit in the hope that Izzy and Anna can settle their differences.
ITV2|1464005700|Coronation Street|||0|0|Soap,Melodrama|Nick is undecided about whether he can cope with moving to Devon and Izzy's revelation that she has been charged with possession of cannabis and assaulting a police officer causes amazement. Elsewhere, Jenny continues to play games with Johnny following her sewing lesson.
ITV2|1464007500|The Ellen DeGeneres Show|||0|0|Talk Show|Actor Ryan Gosling chats about his new film The Nice Guys, which also stars Russell Crowe.
ITV2|1464010800|The Jeremy Kyle Show|23/05/2016 - 1||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.
ITV2|1464015000|The Jeremy Kyle Show|23/05/2016 - 2||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.
ITV2|1464019200|Britain's Got Talent|Live Semi-Final||10|8|General Show,Game Show|Ant and Dec host the first semi-final of this year's contest. The audition process is complete, and has left judges Amanda Holden, David Walliams, Simon Cowell and Alesha Dickson with 45 acts to pick and choose from. Tonight, nine of them will be performing live in the hope of impressing both the panel and the TV audience. The winner of tonight's viewers' vote will automatically go through to the live grand final, before the two runners up face the judges to decide which of them will also win a place.
ITV2|1464024600|Britain's Got Talent Results|Live Results||10|1|General Show,Game Show|Ant and Dec announce the results of tonight's viewers' vote to decide which act will make it through to the grand final. Judges Simon Cowell, David Walliams, Alesha Dixon and Amanda Holden will then select one of the runners up to join them. The show also features a performance by the cast of West End musical Motown.
ITV2|1464026400|You've Been Framed|You've Been Framed! Bounces Back!||0|0|General Show,Game Show|Harry Hill narrates another 60-minute special edition of the comical clip show, applying his unique brand of silly, satirical commentary to a selection of hilarious hi-jinks captured on video by viewers at home.
ITV2|1464030000|Two and a Half Men|Carpet Burns and a Bite Mark||3|3|Sitcom|Charlie is curious about Alan's mysterious love life - until he finds out his brother has been seeing his former wife Judith. He later admits to Rose that he is scared he will miss Jake if the couple patch up their differences and start again. Comedy, starring Charlie Sheen and Jon Cryer.
ITV2|1464031800|Two and a Half Men|Your Dismissive Attitude Toward Boobs||3|4|Sitcom|Berta temporarily moves into the beach house with Charlie and Alan, causing tension to arise between the two men, leading Alan to find his own apartment. Starring Charlie Sheen, Jon Cryer and Conchata Ferrell.
ITV2|1464033600|Family Guy|An App a Day||14|13|Animated Movie,Drama|Peter's newly acquired enthusiasm for smartphone apps inadvertently causes his son Chris to be labelled a sex offender and sent on a rehab course.
ITV2|1464035400|Family Guy|Meet the Quagmires||5|18|Animated Movie,Drama|Death grants Peter his wish to go back in time to 1984, but only for one night. Breaking a date with Lois, he decides to socialise with a famous film star. On his return to the present, he discovers his changes to the timeline have had shocking repercussions.
ITV2|1464037200|Britain's Got More Talent|||10|8|General Show,Game Show|Stephen Mulhern goes behind the scenes of the talent competition's second live semi-final, featuring exclusive chats with celebrity guests, contestants and the judges.
ITV2|1464040800|Family Guy|Airport '07||5|12|Animated Movie,Drama|Quagmire loses his job as a pilot and has trouble finding alternative employment, so Peter and Cleveland hatch a plan to get him reinstated - which entails jeopardising an airliner full of passengers. With the guest voice of Hugh Hefner.
ITV2|1464042600|American Dad|A Jones for a Smith||6|11|Animated Movie,Drama|Stan complains that liberal social programmes are a waste of money and criticises Francine for helping at the local homeless shelter - until he develops a crack cocaine addiction and suddenly has a change of heart.
ITV2|1464044100|American Dad|May the Best Stan Win||6|12|Animated Movie,Drama|Francine is swept off her feet by a romantic cyborg version of her husband who has come back from the future, and the encounter forces her to question her relationship with the real Stan. Meanwhile, Roger directs Steve and his friends in a remake of cult classic adventure movie The Goonies.
ITV2|1464045900|The Cleveland Show|The Hurricane||3|2|Animated Movie,Drama|The Brown and Tubbs families try to salvage what is left of their holidays when a storm hits Stoolbend, while Cleveland Jr makes a surprising announcement about his religious beliefs.(n)
ITV2|1464047700|The Cleveland Show|A Nightmare on Grace Street||3|3|Animated Movie,Drama|Cleveland and Rallo worry they might be cowards after they are both sent home from sleepovers for getting scared. Donna decides to tackle the issue by taking them to spend the night at a haunted house, where she hopes to prove they are both braver than they think. Meanwhile, Roberta is trapped in a love triangle between a vampire and a werewolf.(n)
ITV2|1464049200|Celebrity Juice|||15|10|Comedy|Funnyman Jimmy Carr and Bang on the Money presenting duo Rickie Haywood-Williams and Melvin Odoom join in the fun, with Holly Willoughby, Fearne Cotton and Gino D'Acampo.(n)
ITV2|1464051900|@elevenish|||1|10|Comedy|Topical comedy series in which a cast of stand-ups, character actors and comedy groups share their thoughts on the past seven days through monologues, sketches and commentary.(n)
ITV2|1464053400|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.(n)
ITV2|1464066000|The Hot Desk|The Hot Desk: Adam Lambert||0|0|General Music,Ballet,Dance|Exclusive interviews with the hottest names in music and entertainment. Behind the desk today is US singer, songwriter and stage actor Adam Lambert.(n)
ITV2|1464066600|Dinner Date|Martin||1|30|Cooking|Londoner Martin picks three blind dates from five potential partners, based entirely on the menus they have created. When the three dinners have been eaten, he decides who he wants to see again. Narrated by Charlotte Hudson.(n)
ITV2|1464069600|The Ellen DeGeneres Show|||0|0|Talk Show|Actor Ryan Gosling chats about his new film The Nice Guys, which also stars Russell Crowe.(n)
ITV2|1464072600|Emmerdale|||0|0|Soap,Melodrama|Lawrence demands that Ronnie leave his family alone, only to find the plumber knows things he would rather keep secret. Doug tries to give Laurel a break from her worries, and Chrissie is delighted when her divorce comes through. Vanessa is less than thrilled when Carly invites Tracy to come and live with them, and Sam fears Megan is considering giving Jai another chance.(n)
ITV2|1464074400|Coronation Street|||0|0|Soap,Melodrama|Long-running drama with the residents of England's most famous cobbled street.(n)
ITV2|1464076200|Coronation Street|||0|0|Soap,Melodrama|With Johnny nowhere to be found, Roy offers to walk Carla down the aisle, but as she comes face to face with the groom, the bride tells Nick she wants to speak to him in private. Will the ceremony go ahead?.(n)
ITV2|1464078000|Psych|Black and Tan: A Crime of Fashion||2|15|Comedy|Shawn and Gus are plunged into the world of fashion as they investigate the murder of a designer. Detective comedy, starring James Roday and Dule Hill.(n)
ITV2|1464081000|Britain's Got Talent|Live Semi-final Two||10|9|General Show,Game Show|Ant and Dec present the second live semi-final, as nine more of the 45 chosen acts compete to impress judges Amanda Holden, David Walliams, Simon Cowell and Alesha Dixon and secure the all-important viewers' vote. At stake is the chance to appear at this year's Royal Variety Performance and win a life-changing cash prize of £250,000, with the act with the highest public vote going through automatically, while two runners-up fight it out for the judges' favour.(n)
ITV2|1464086700|Britain's Got Talent Results|||10|2|General Show,Game Show|Ant and Dec announce the act with the highest number of public votes, automatically going through to the final. Simon Cowell, David Walliams, Amanda Holden and Alesha Dixon then decide which of the contestants in second and third place they want to see again. Plus, American pop-rock band One Republic perform.(n)
ITV2|1464088500|Emmerdale|||0|0|Soap,Melodrama|Lawrence demands that Ronnie leave his family alone, only to find the plumber knows things he would rather keep secret. Doug tries to give Laurel a break from her worries, and Chrissie is delighted when her divorce comes through. Vanessa is less than thrilled when Carly invites Tracy to come and live with them, and Sam fears Megan is considering giving Jai another chance.(n)
ITV2|1464090300|Coronation Street|||0|0|Soap,Melodrama|Long-running drama with the residents of England's most famous cobbled street.(n)
ITV2|1464092100|Coronation Street|||0|0|Soap,Melodrama|With Johnny nowhere to be found, Roy offers to walk Carla down the aisle, but as she comes face to face with the groom, the bride tells Nick she wants to speak to him in private. Will the ceremony go ahead?.(n)
ITV2|1464093900|The Ellen DeGeneres Show|24/05/2016||0|0|Talk Show|The comedienne is joined in the studio by Christina Aguilera, currently a coach on the US version of The Voice, along with Pete's Dragon star Bryce Dallas Howard and beauty expert Kym Douglas.(n)
ITV2|1464097200|The Jeremy Kyle Show|24/05/2016 - 1||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.(n)
ITV2|1464101400|The Jeremy Kyle Show|24/05/2016 - 2||0|0|Talk Show|The host invites guests to air their differences over family and relationship issues, and provides them with his own brand of no-nonsense advice.(n)
ITV2|1464105600|Britain's Got Talent|Live Semi-final Two||10|9|General Show,Game Show|Ant and Dec present the second live semi-final, as nine more of the 45 chosen acts compete to impress judges Amanda Holden, David Walliams, Simon Cowell and Alesha Dixon and secure the all-important viewers' vote. At stake is the chance to appear at this year's Royal Variety Performance and win a life-changing cash prize of £250,000, with the act with the highest public vote going through automatically, while two runners-up fight it out for the judges' favour.(n)
ITV2|1464111000|Britain's Got Talent Results|||10|2|General Show,Game Show|Ant and Dec announce the act with the highest number of public votes, automatically going through to the final. Simon Cowell, David Walliams, Amanda Holden and Alesha Dixon then decide which of the contestants in second and third place they want to see again. Plus, American pop-rock band One Republic perform.(n)
ITV2|1464112800|You've Been Framed|||28|13|General Show,Game Show|Harry Hill narrates another selection of comical home videos, provided by viewers armed with everything from drones to selfie-sticks. Among tonight's highlights are a man falling off a bridge into a canal, a lion jumping into a car during a safari, and a student who finds an unwelcome surprise in her toilet.(n)
ITV2|1464114600|You've Been Framed|||28|2|General Show,Game Show|Harry Hill narrates another selection of comical mishaps filmed by viewers, including an unusual take on Ninja Warrior UK, a preview of what Ant and Dec might look like in their sixties, and a fine example of why riding a bicycle is not the best time to take a selfie. Plus, a family is soaked by what appears to be an exploding colon.(n)
ITV2|1464116400|Two and a Half Men|We Called It Mr Pinky||3|5|Sitcom|Rose tells Charlie he is unable to sustain a lasting relationship with a woman because of his attitude to his mother, and Jake seeks advice about a girl at school. Starring Charlie Sheen, Jon Cryer and Angus T Jones.(n)
ITV2|1464118200|Two and a Half Men|Hi, Mr Horned One||3|6|Sitcom|Charlie continues to date an attractive Satan worshipper - despite Alan's warnings - but when she threatens to put a curse on his manhood, he begins to see sense. Starring Charlie Sheen, Jon Cryer and Jodi Lyn O'Keefe.(n)
ITV2|1464120000|Family Guy|The Simpsons Guy - Part One||13|1|Animated Movie,Drama|The Griffin family find themselves stuck in Springfield, home to The Simpsons, after fleeing Quahog when Peter faces a backlash over a misogynistic comic strip.(n)
ITV2|1464121800|Family Guy|The Simpsons Guy - Part Two||13|1|Animated Movie,Drama|Conclusion of the story in which the Griffin family are stuck in Springfield, home to The Simpsons, after Peter creates a controversial comic strip.(n)
ITV2|1464123600|Britain's Got More Talent|||0|0|General Show,Game Show|Stephen Mulhern covers the reactions, gossip from the judges, and behind the scenes drama as the live semi-finals continue.(n)
ITV2|1464127200|Family Guy|Baking Bad||13|3|Animated Movie,Drama|Peter and Lois go into business together, opening a cookie store. However, tensions rise when Peter devises his own way of attracting more customers. Adult animation, featuring the voices of Seth MacFarlane and Alex Borstein.(n)
ITV2|1464129000|Family Guy|Bill and Peter's Bogus Journey||5|13|Animated Movie,Drama|Peter is upset to learn that Lois has slept with his new friend Bill Clinton and decides to retaliate by having an affair of his own - but soon realises he loves her too much to ever be unfaithful. Meanwhile, Lois and Stewie try to potty-train Brian.(n)
ITV3|1463871600|Trial & Retribution|Ghost Train - Part One||12|3|Detective,Thriller|Part one of two. A girl falls to her death from a Ferris wheel in what appears to be a tragic accident, but a fortune-teller from the funfair reveals she suspects foul play. DS Satchell is embarrassed to discover the woman is a distant relative and finds himself working alone to prove a murder has been committed - until a second death confirms his suspicions. Jane Lapotaire guest stars.
ITV3|1463875500|Northern Lights|||1|3|General Movie,Drama|The feuding brothers-in-law attend a school reunion, where things almost turn nasty as Colin has a run-in with an enemy from his childhood. Meanwhile, Howie bumps into an old flame and quickly rekindles their former relationship - jeopardising his marriage in the process. It's up to his oldest mate to decide whether to dish the dirt to Pauline and betray his friend's trust. Comedy drama, starring Robson Green.
ITV3|1463878800|ITV3 Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV3|1463880600|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.
ITV3|1463893200|On the Buses|The New Nurse||5|8|Sitcom|The new depot nurse moves in as the Butlers' lodger - causing problems for Arthur. Vintage comedy, starring Reg Varney and Michael Robbins.
ITV3|1463894700|The Return of Sherlock Holmes|The Empty House||1|1|Mystery|The great detective reveals to a startled Watson how he defeated Moriarty and cheated death beneath the waters of the Reichenbach Falls. Period drama, marking Edward Hardwicke's debut as Holmes' indefatigable chronicler.
ITV3|1463898000|Heartbeat|Scent of a Kill||13|14|General Movie,Drama|Dr Merrick faces a testing time when a terrified hospital patient claims her husband is trying to kill her, but Merton seems reluctant to get involved, while Vernon picks up a bargain all-purpose pest-control solution, enlisting David's help in his eradication mission. Gina's cousin Diane arrives to help her and Phil with the wedding preparations - much to the delight of PC Crane, who is instantly smitten. Rural drama, starring Aislin McGuckin, Tricia Penrose and Mark Jordon.
ITV3|1463901900|Heartbeat|Daniel||13|15|General Movie,Drama|Steve is forced to cover for Phil when the father-to-be discovers Gina has gone into labour two months early and rushes to the hospital to help with the nerve-racking delivery. Meanwhile, Merton is excited when it appears a drug dealer could soon be brought to justice. Drama, starring Mark Jordon, Tricia Penrose and Duncan Bell.
ITV3|1463905800|Inspector Morse|The Wolvercote Tongue||2|1|Detective,Thriller|An American tourist's body is discovered in her hotel room, apparently dead from a heart attack - but a valuable Anglo-Saxon jewel she intended to donate to the Ashmolean Museum is missing and several interested parties are acting strangely. John Thaw and Kevin Whately star, with Simon Callow, Roberta Taylor and Kenneth Cranham.
ITV3|1463913900|Foyle's War|They Fought in the Fields||3|3|Detective,Thriller|A farmer's murder and the crash landing of an enemy plane lead Foyle to investigate the activities of a group of land girls, and the detective begins to suspect the captured German airmen have something to hide. Stella Gonet and James Wilby guest star in the wartime drama, with Michael Kitchen, Anthony Howell and Honeysuckle Weeks.
ITV3|1463921400|Columbo: Any Old Port in a Storm||1973|0|0|Police,Crime Drama|A vineyard owner's financial security is jeopardised when his playboy younger brother threatens to sell the family winery. He resorts to killing his sibling and rigging the death scene to look like a scuba-diving accident. However, the crumpled cop sees through the ruse and in the process reveals he is something of a wine buff himself. Detective drama, with Peter Falk, Donald Pleasence and Julie Harris.
ITV3|1463928600|Agatha Christie's Marple|Towards Zero||3|4|Mystery|A gathering at the Devon estate of Miss Marple's old school friend Lady Tressilian leads to murder when the eccentric Mr Treves tells the story of an unconvicted child killer. Miss Marple is on hand to assist Supt Mallard of the local constabulary, but not before a second victim is claimed. Mystery, starring Geraldine McEwan, with guest appearances by Eileen Atkins, Tom Baker, Paul Nicholls, Alan Davies and Greg Wise, with a cameo by former British number-one tennis player Greg Rusedski.
ITV3|1463936100|Margery and Gladys|||0|0|Comedy|Two mismatched elderly ladies interrupt a burglary and hit the culprit over the head in a panic, leaving him for dead before going on the run. As they head for Blackpool, a series of unexpected developments soon make things worse - and then there's the police, who are hot on their heels. One-off comedy, starring Penelope Keith, June Brown, Alan David and Marcia Warren.
ITV3|1463943600|Rosemary & Thyme|The Memory of Water||2|0|Mystery|The amateur sleuths are hired to bring a mansion's walled garden back to life, with help from inmates of the local prison. Events take a sinister turn when the owner's cousin is found drowned in the local fast-flowing river - and become even more mysterious when, just before the inquest, Rosemary sees the dead man alive. Feature-length edition of the mystery drama, starring Felicity Kendal and Pam Ferris.
ITV3|1463950800|Ghostboat|||1|2|General Movie,Drama|Concluding part. Hardy finds himself fighting to stop events as the forgotten happenings of 1943 start to have deadly consequences. Struggling to hang on to their identities, the Scorpion's latter-day crew discover that what is waiting for them under the grey waters of the Baltic Sea is far worse than the Russian submarines they expected. Drama, with David Jason, Ian Puleston-Davies and Tony Haygarth.
ITV3|1463956500|Agatha Christie's Marple|Towards Zero||3|4|Mystery|A gathering at the Devon estate of Miss Marple's old school friend Lady Tressilian leads to murder when the eccentric Mr Treves tells the story of an unconvicted child killer. Miss Marple is on hand to assist Supt Mallard of the local constabulary, but not before a second victim is claimed. Mystery, starring Geraldine McEwan, with guest appearances by Eileen Atkins, Tom Baker, Paul Nicholls, Alan Davies and Greg Wise, with a cameo by former British number-one tennis player Greg Rusedski.
ITV3|1463963700|Blue Murder|Having It All||5|1|Detective,Thriller|DCI Janine Lewis struggles to balance family life with an investigation into the murder of a cheerleading coach. Initial suspicion falls on the victim's husband, whose bloodied clothes are found near the crime scene, but the discovery of an affair suggests someone else may have had a motive. Guest starring Coronation Street's Chris Gascoyne.
ITV3|1463966700|May the Best House Win|South Yorkshire and Derbyshire||5|12|Game Show,Quiz|The competition heads to South Yorkshire and Derbyshire, where glamorous gran Liz Treece, model-agency owner Jo Webster, renewable energy fanatic Mark Woodward and singleton Nigel Fox score one another's properties. They open their doors to a modern detached home, a renovated chapel, a converted barn and farmhouse, and a bachelor pad, in the hope of winning the £1,000 prize. Narrated by Guy Porritt.
ITV3|1463970000|May the Best House Win|Cambridgeshire & Suffolk 2||5|19|Game Show,Quiz|Four homeowners in Cambridgeshire and Suffolk rate one another's houses in a bid to win £1,000. The homes under inspection are Claire Avenal's heart-filled terraced property in Newmarket, Katie Lancashire's modern detached house, landlord David Utting's pub and Aletta Wilson's spacious abode, converted from a former Salvation Army church hall. Narrated by Guy Porritt.
ITV3|1463973000|On the Buses|Lost Property||5|9|Sitcom|A woman arrives at the depot to claim her lost property, but Stan and Jack have already eaten it. Comedy, starring Reg Varney and Bob Grant.
ITV3|1463974500|On the Buses|Stan's Uniform||5|10|Sitcom|Stan gets a new uniform and is proud to wear it - until he sits on a freshly painted chair. Classic comedy, starring Reg Varney.
ITV3|1463976000|Judge Judy|22/05/2016 - 1||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.
ITV3|1463977500|Judge Judy|22/05/2016 - 2||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.
ITV3|1463978700|ITV3 Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV3|1463979600|In Loving Memory|Gone Dancing||1|3|Comedy|Ivy has hopes for nephew Billy's chances with the girls at the local dance. Comedy set in an undertakers, starring Thora Hird.
ITV3|1463981100|Heartbeat|Oscar's Birthday||17|24|General Movie,Drama|Two new residents put PC Mason in an awkward position both professionally and personally and, while the village rallies round to celebrate Blaketon's birthday, he gets more than he expected when Gina goes into labour. David decides to learn to play the piano. Rural police drama set in the rustic backwater of Aidensfield, Yorkshire. Starring Joe McFadden, Tricia Penrose and Derek Fowlds.
ITV3|1463985000|Where the Heart Is|The Games We Play||8|4|General Movie,Drama|Anna is unsure whether she should tell Luke the truth about his chances of recovery after his near-fatal rugby accident, and Ozias Harding's persistent bullying forces Billy to resign from the factory, leading Nathan to take revenge against the businessman by asking out his daughter Alice. Lesley Dunlop, Brian Capron and Andrew Paul star.
ITV3|1463988600|The Royal|These Foolish Things||8|3|General Movie,Drama|Weatherill treats a schoolgirl whose crush on a teacher has spiralled out of control, while Ormerod and Ellis launch a daring cliff rescue when a family picnic goes awry. Jack and Alun use a map to hunt for buried treasure underneath the hospital, and an old friend of Matron is taken ill. Sixties-set medical drama, starring Amy Robbins, Robert Daws, Neil McDermott and Wendy Craig.
ITV3|1463992500|Judge Judy|23/05/2016 - 1||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.
ITV3|1463994000|Judge Judy|23/05/2016 - 2||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.
ITV3|1463995500|Judge Judy|23/05/2016 - 3||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.
ITV3|1463997300|Murder, She Wrote|Benedict Arnold Slipped Here||4|18|Mystery|Cabot Cove becomes the scene of deadly competition when an eccentric recluse dies, and Jessica is given the dubious honour of executing the woman's will. Starring Angela Lansbury.
ITV3|1464000900|The Return of Sherlock Holmes|The Abbey Grange||1|2|Mystery|Captain Jack Crocker, a robust seafaring man, is implicated in the murder of beautiful aristocrat Lady Brackenstall's abusive husband. Drama, guest starring Oliver Tobias, with Jeremy Brett, Edward Hardwicke and Anne Louise Lambert.
ITV3|1464004800|Heartbeat|Family Matters||18|1|General Movie,Drama|An encounter with a gang of armed men presents Miller with a difficult dilemma that puts his professional and personal future in jeopardy. Mason and Wetherby struggle to deal with student protesters who are furious at the presence of a suspected Nazi collaborator in the town, and the situation escalates further when an attempt is made on the man's life. John Duttine and Joe McFadden star.
ITV3|1464008700|The Royal|Any Old Iron||8|4|General Movie,Drama|Continuing the final series of the hospital drama after a two-year break. Susie Dixon's head is turned by a rich playboy, with devastating consequences for Mrs Middleditch when the negligent nurse administers the wrong blood during a transfusion. Ormerod is called out by the coastguard to rescue a grieving widow who has got into difficulty on her yacht, and Jack and Alun find themselves looking after a horse after it tramples its owner. Robert Daws, Sarah Beck Mather, Susan Hampshire and Gareth Hale star.
ITV3|1464012300|Where the Heart Is|Little Boy Blue||8|5|General Movie,Drama|Luke arrives back home in a wheelchair, but quickly becomes frustrated and takes his anger out on David. Charlie tries to avoid his daughter Charlotte when she returns from Italy and Nathan convinces Alice to keep their relationship secret - a move which drives her to accept a date with Joe.
ITV3|1464016200|In Loving Memory|The Rivals||1|4|Comedy|Ivy is distraught to find that a rival undertaker is setting up in town. Comedy, starring Thora Hird.
ITV3|1464018600|On the Buses|A Thin Time||5|14|Sitcom|Beryl describes her ideal man, leaving Arthur dejected because he does not even begin to measure up. Reg Varney stars.
ITV3|1464020400|George and Mildred|Days of Beer and Rosie||4|2|Sitcom|The thought of being a step-grandmother leaves Mildred distraught. Comedy, starring Brian Murphy and Yootha Joyce.
ITV3|1464022500|Heartbeat|Family Matters||18|1|General Movie,Drama|An encounter with a gang of armed men presents Miller with a difficult dilemma that puts his professional and personal future in jeopardy. Mason and Wetherby struggle to deal with student protesters who are furious at the presence of a suspected Nazi collaborator in the town, and the situation escalates further when an attempt is made on the man's life. John Duttine and Joe McFadden star.
ITV3|1464026400|Murder, She Wrote|Just Another Fish Story||4|19|Mystery|Jessica invests in an upmarket New York seafood restaurant, but unfortunately the maitre d' is murdered shortly afterwards, leaving her facing the double dilemma of recouping her cash outlay and catching the killer. Guest starring Sonny Bono and Brenda Vaccaro.
ITV3|1464030000|Lewis|Entry Wounds||0|0|Detective,Thriller|The last run of the detective drama ended with Lewis (Kevin Whately) starting a new life away from the force, but it seems that peace and quiet doesn't suit him - which is just as well, as newly promoted DI Hathaway (Laurence Fox) is struggling to find a sidekick, and within just four weeks is already on to his second sergeant, DS Lizzie Maddox (Angela Griffin). So, Chief Superintendent Innocent (Rebecca Front) decides to reunite the former partners to look into the murder of a neurosurgeon, a case with potential links to the worlds of animal rights and blood sports. Suspicion falls on glamorous widow Erica (Kara Tointon), but it turns out there are plenty of other people in the victim's inner circle who were driven by fear and loathing.
ITV3|1464037200|Wycliffe|Time Out||5|2|Detective,Thriller|A prostitute's client confesses to the murder of another working girl before vanishing into the night, leaving Wycliffe with the tricky task of tracking him down before he kills again. Detective drama, starring Jack Shepherd.
ITV3|1464040800|The Knock|||2|6|General Movie,Drama|The net begins to close on Webster as Bill flies to Portugal to take a closer look at his operation, while by the team carry out a raid on Rufus Teague.
ITV3|1464045300|Cold Blood|||0|0|General Movie,Drama|Matthew Kelly stars as a serial killer who has spent his 15 years in prison playing a game of psychological cat-and-mouse with his captors. One of Britain's most notorious murderers, Brian Wicklow is vilified by the Press and despised by fellow inmates - not least because detectives have never found the body of his last victim. But then, out of the blue, he decides he wants to talk to the police. John Hannah, Jemma Redgrave and David Calder co-star.(n)
ITV3|1464049800|On the Buses|Bye Bye Blakey||6|6|Sitcom|Stan and Jack eavesdrop on Blakey's medical - and completely misinterpret its findings. Comedy, starring Reg Varney, Bob Grant and Stephen Lewis.(n)
ITV3|1464051600|ITV3 Nightscreen|||0|0|General Education,Science|Text-based information service.(n)
ITV3|1464053400|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.(n)
ITV3|1464066000|In Loving Memory|The Rivals||1|4|Comedy|Ivy is distraught to find that a rival undertaker is setting up in town. Comedy, starring Thora Hird.(n)
ITV3|1464067500|Heartbeat|Family Matters||18|1|General Movie,Drama|An encounter with a gang of armed men presents Miller with a difficult dilemma that puts his professional and personal future in jeopardy. Mason and Wetherby struggle to deal with student protesters who are furious at the presence of a suspected Nazi collaborator in the town, and the situation escalates further when an attempt is made on the man's life. John Duttine and Joe McFadden star.(n)
ITV3|1464071400|Where the Heart Is|Little Boy Blue||8|5|General Movie,Drama|Luke arrives back home in a wheelchair, but quickly becomes frustrated and takes his anger out on David. Charlie tries to avoid his daughter Charlotte when she returns from Italy and Nathan convinces Alice to keep their relationship secret - a move which drives her to accept a date with Joe.(n)
ITV3|1464075000|The Royal|Any Old Iron||8|4|General Movie,Drama|Continuing the final series of the hospital drama after a two-year break. Susie Dixon's head is turned by a rich playboy, with devastating consequences for Mrs Middleditch when the negligent nurse administers the wrong blood during a transfusion. Ormerod is called out by the coastguard to rescue a grieving widow who has got into difficulty on her yacht, and Jack and Alun find themselves looking after a horse after it tramples its owner. Robert Daws, Sarah Beck Mather, Susan Hampshire and Gareth Hale star.(n)
ITV3|1464078900|Judge Judy|24/05/2016 - 1||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.(n)
ITV3|1464080400|Judge Judy|24/05/2016 - 2||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.(n)
ITV3|1464081900|Judge Judy|24/05/2016 - 3||0|0|General Education,Science|Real-life small-claims cases on issues affecting family life, presided over by outspoken former New York judge Judy Sheindlin.(n)
ITV3|1464083700|Murder, She Wrote|Just Another Fish Story||4|19|Mystery|Jessica invests in an upmarket New York seafood restaurant, but unfortunately the maitre d' is murdered shortly afterwards, leaving her facing the double dilemma of recouping her cash outlay and catching the killer. Guest starring Sonny Bono and Brenda Vaccaro.(n)
ITV3|1464087300|The Return of Sherlock Holmes|The Man with the Twisted Lip||1|5|Mystery|A woman asks Holmes to search for her missing husband, a businessman who was last seen peering from the window of an opium den in London's notorious Limehouse area. Suspicion falls on a well-known local beggar - but his innocence is eventually proved in bizarre fashion. Period drama, starring Jeremy Brett.(n)
ITV3|1464091500|Heartbeat|England Expects||18|2|General Movie,Drama|A notorious burglar escapes from prison and returns to Aidensfield to pursue a vendetta against Ashfordly police. Roping in two local boys, the villain dupes them into helping him carry out his plan while PC Mason desperately tries to find him before he strikes again. Dawn sets Joyce up on a date with PC Younger - but is oblivious to the fact that the young copper actually has feelings for her. George Cole guest stars, with Joe McFadden and John Duttine.(n)
ITV3|1464095100|The Royal|Should I Stay or Should I Go Now||8|5|General Movie,Drama|Timid new student nurse Faye Clark is faced with a trying first day when a model collapses after taking magic mushrooms. Lizzie falls for an injured motorcycle stuntman who is convinced he is destined to live fast and die young due to a hereditary condition - but Ormerod comes up with a different diagnosis. Lauren Drummond, Michelle Hardwick, James Daffern and Robert Daws star.(n)
ITV3|1464099000|Where the Heart Is|Skin Deep||8|6|General Movie,Drama|A patient's wife accuses Sally of having an affair with her husband, putting pressure on the nurse's career and marriage, while Nathan and Joe find out the truth about Alice's two-timing and a bored Alan discovers he has won the star prize on a scratch card. Ex-EastEnder Martin Kemp guest stars.(n)
ITV3|1464102900|In Loving Memory|Pork||1|5|Comedy|Ivy attends the funeral of a friend's husband who had an unfortunate incident with a tram. Comedy, starring Thora Hird.(n)
ITV3|1464105000|On the Buses|The New Telly||5|12|Sitcom|Stan splashes out on a new colour television for the family, but has problems disposing of the old one. Vintage comedy, starring Reg Varney.(n)
ITV3|1464106800|George and Mildred|You Must Have Showers||4|3|Sitcom|Mrs Roper wants to install a shower, but a lack of cash forces a compromise on costs - and workmanship. Brian Murphy and Yootha Joyce star.(n)
ITV3|1464108900|Heartbeat|England Expects||18|2|General Movie,Drama|A notorious burglar escapes from prison and returns to Aidensfield to pursue a vendetta against Ashfordly police. Roping in two local boys, the villain dupes them into helping him carry out his plan while PC Mason desperately tries to find him before he strikes again. Dawn sets Joyce up on a date with PC Younger - but is oblivious to the fact that the young copper actually has feelings for her. George Cole guest stars, with Joe McFadden and John Duttine.(n)
ITV3|1464112800|Murder, She Wrote|Showdown in Saskatchewan||4|20|Mystery|Jessica investigates a mysterious death, the repercussions of which are causing unrest among the riders at a rodeo. Starring Angela Lansbury, Kristy McNichol and Larry Wilcox.(n)
ITV3|1464116400|Lewis|The Lions of Nemea||8|0|Detective,Thriller|Hathaway appears to have got over his fear of Lewis treading over his newly promoted toes. Their opposites have attracted in the past, and there seems no reason to suspect that they won't now the younger man has got used to the idea of his former mentor coming out of retirement to lend him a hand. Even DS Maddox isn't getting on Hathaway's nerves quite as much, so this rejuvenated trio sets out to discover who murdered American classics student Rose Anderson, whose body has been hauled from the canal with neck and abdomen wounds. Nevertheless, a few red herrings threaten to get in their way of landing the killer. Kevin Whately, Laurence Fox and Angela Griffin star.(n)
ITV3|1464123600|Wycliffe|Standing Stone||5|3|Detective,Thriller|Sophie, the wife of one of Kersey's friends, goes missing after an evening class and soon her tutor is found murdered. The detectives step in to investigate but the clues lead to standing stones linked to the entrance to hell in local superstition. Jack Shepherd and Helen Masters star.(n)
ITV3|1464127200|The Knock|||2|7|General Movie,Drama|Barry refuses to accept that his relationship with Diane is over, Katherine feels humiliated by the outcome of the Short case, and Webster infuriates his partners in crime.(n)
ITV4|1463871600|FYI Daily|21/05/2016 - 4||0|0|News Magazine,Current Affairs|
ITV4|1463871900|State of Play||2009|0|0|Detective,Thriller|A hard-nosed journalist investigating the murder of a congressman's intern discovers a connection between the tragedy and the death of a petty crook on the same evening. As he works to get to the bottom of the story, the reporter uncovers a political conspiracy that places him in a precarious and potentially life-threatening position. Thriller, starring Russell Crowe, Ben Affleck, Helen Mirren and Rachel McAdams.
ITV4|1463876100|Hell on Wheels|Blood Moon||2|9|Western|Part one of two. The townsfolk celebrate the completion of the bridge. Meanwhile Cullen suspects the Sioux are preparing to attack and Durant has a deadly task for Elam.
ITV4|1463879400|Ax Men|The Mouth from the South||4|15|Documentary|Conflict between Craig and Dave at Rygaard threatens to tear the crew apart, and at Papac Alaska, Joe and Coatsy get a chance to make amends.
ITV4|1463882400|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.
ITV4|1463893200|Football's Greatest: Thierry Henry|||0|0|General Sports|A profile of the former striker, who won a number of honours with France, Arsenal and Barcelona.
ITV4|1463893500|Motorway Patrol|||0|0|Documentary|Documentary following members of the New Zealand highway patrol as they witness the best and worst behaviour on the nation's busiest motorway.
ITV4|1463895300|Fifth Gear|||26|6|Motoring|The team investigates car culture in Romania, testing extreme off-road vehicles in its countryside and ski resorts and meeting a classic car restorer in Bucharest.
ITV4|1463898900|Fifth Gear|||26|1|Motoring|Tiff Needell and Vicki Butler-Henderson take part in a unique car versus plane challenge as Red Bull Air Race champion Nigel Lamb takes on a Lamborghini Aventador. The plane is clearly faster, but there is the small matter of cornering. On the track, the VW Golf R is put up against the Subaru WRX STi to see which is faster. Plus, Jonny Smith becomes an official test driver for the day and the team tests Citroen's tiny C1 city car.
ITV4|1463902500|Pawn Stars|Every Day I'm Shufflin'||8|25|General Show,Game Show|An official film prop from The Godfather makes its way into the shop, as does a piece of 1950s bowling equipment. Meanwhile, tensions build between Chumlee and the Old Man. Reality programme chronicling the daily activities at the World Famous Gold & Silver Pawn Shop in Las Vegas.
ITV4|1463904000|Pawn Stars|The Bald and the Beautiful||8|0|General Show,Game Show|A coat custom-made for Elvis Presley makes for an excited team. Plus, Chumlee gives a Mercedes Benz golf cart the once over. Reality programme chronicling the daily activities at the World Famous Gold & Silver Pawn Shop in Las Vegas.
ITV4|1463905800|Live French Open Tennis|2016 Day One||0|0|Tennis|John Inverdale presents coverage of the opening day of the second Grand Slam event of the year, staged at Roland Garros in Paris, featuring first-round matches from both the men's and women's draws. The opening round of last year's tournament saw a number of seeded players eliminated at the first time of asking, with Grigor Dimitrov among five players to lose in the men's draw, and Eugenie Bouchard one of six ladies to suffer an early exit. With analysis from Marion Bartoli, Jim Courier, Mark Petchey, Fabrice Santoro and Sam Smith, commentary by Nick Mullins and reports from Celina Hinchcliffe.
ITV4|1463947200|Premiership Rugby Union|2015/16 Semi-Finals||0|0|Rugby Union - Domestic|Mark Durden-Smith and David Flatman present highlights of the semi-finals, which were Saracens v Leicester Tigers at Allianz Park and Exeter Chiefs v Wasps at Sandy Park.
ITV4|1463950800|Raw Deal||1986|0|0|Detective,Thriller|An FBI agent is discharged for insubordination after assaulting a suspect, and ends up reduced to being the sheriff of a backwater Southern town. He is later offered his old job back - on the condition he will infiltrate a gang of Chicago mobsters and bring their leader to justice for killing the son of the Bureau's chief. Action thriller, with Arnold Schwarzenegger, Sam Wanamaker, Kathryn Harrold, Ed Lauter and Darren McGavin.
ITV4|1463954400|FYI Daily|22/05/2016 - 1||0|0|News Magazine,Current Affairs|
ITV4|1463954700|Raw Deal||1986|0|0|Detective,Thriller|An FBI agent is discharged for insubordination after assaulting a suspect, and ends up reduced to being the sheriff of a backwater Southern town. He is later offered his old job back - on the condition he will infiltrate a gang of Chicago mobsters and bring their leader to justice for killing the son of the Bureau's chief. Action thriller, with Arnold Schwarzenegger, Sam Wanamaker, Kathryn Harrold, Ed Lauter and Darren McGavin.
ITV4|1463958600|Red Heat||1988|0|0|Adventure|A Russian detective travels to America to oversee the extradition of a Georgian drug baron responsible for supplying cocaine in Moscow. He is teamed up with a hostile Chicago cop, but when their prisoner kills an officer and escapes, they put aside their mutual mistrust to bring him to justice. Action thriller, starring Arnold Schwarzenegger, James Belushi, Peter Boyle, Laurence Fishburne and Ed O'Ross.
ITV4|1463962200|FYI Daily|22/05/2016 - 2||0|0|News Magazine,Current Affairs|
ITV4|1463962500|Red Heat||1988|0|0|Adventure|A Russian detective travels to America to oversee the extradition of a Georgian drug baron responsible for supplying cocaine in Moscow. He is teamed up with a hostile Chicago cop, but when their prisoner kills an officer and escapes, they put aside their mutual mistrust to bring him to justice. Action thriller, starring Arnold Schwarzenegger, James Belushi, Peter Boyle, Laurence Fishburne and Ed O'Ross.
ITV4|1463966400|Tommy Cooper|||1|6|Comedy|Patrick Cargill and Trisha Noble join the incomparable comedian as he performs a variety of sketches.
ITV4|1463968500|ITV4 Nightscreen|||0|0|General Education,Science|Text-based information service.
ITV4|1463968800|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.
ITV4|1463979600|Tommy Cooper|||0|0|Comedy|The comedian performs a variety of sketches and magic tricks.
ITV4|1463981400|Minder|The Dessert Song||1|10|General Movie,Drama|Arthur and Terry rescue Greek-Cypriot Charlie from a beating and learn that his cousin is being threatened by another relative who wants to take over their restaurant. Encouraged by Charlie who is vowing revenge, Terry takes a job in the establishment to try to catch the tormentors red-handed.
ITV4|1463985300|The Chase|23/05/2016||0|0|Quiz Show|Bradley Walsh presents as four contestants pit their wits against ruthless quiz genius the Chaser in the hope of winning a potential prize pot worth thousands of pounds. They work as a team and play strategically to answer general knowledge questions against the clock and race down the game board to the exit without being caught.
ITV4|1463988900|Storage Wars: Texas|Bubbapocalypse Now||2|8|Documentary|The bidders compete over collectible dolls, antiques and a strange coin, which supposedly has the means to prevent the end of the world.
ITV4|1463990400|Storage Wars: Texas|Night of the Pondering Dead||2|9|Documentary|The buyers attend auctions in Ponder, but face stiff competition from the locals, who seem to have inside knowledge on the contents of the lockers.
ITV4|1463992200|Live French Open Tennis|2016 Day Two||0|0|Tennis|John Inverdale presents coverage of day two of the second Grand Slam event of the year, staged at Roland Garros in Paris, featuring the latest matches in the first round. Eventual champions Stan Wawrinka and Serena Williams both recorded straight-sets victories in the opening round of last year's tournament, with Wawrinka defeating Marsel Ilhan 6-3, 6-2, 6-3, and Williams recording a 6-2, 6-3 win over Andrea Hlavackova. With analysis from Marion Bartoli, Jim Courier, Mark Petchey, Fabrice Santoro and Sam Smith, commentary by Nick Mullins and reports from Celina Hinchcliffe.
ITV4|1464033600|MotoGP Highlights|2016 Italian Grand Prix||0|0|Motorcycling|The Italian Grand Prix. Action from the sixth round of the season, which was staged at the Mugello Circuit in Tuscany, Italy.
ITV4|1464037200|Heartbreak Ridge||1986|0|0|Adventure,War|A hellraising US marine sergeant is assigned to whip a squad of raw recruits into shape for the invasion of Grenada in 1983 - but his old-fashioned methods meet with disapproval from superior officers. Action adventure, directed by and starring Clint Eastwood. With Marsha Mason, Everett McGill, Moses Gunn and Bo Svenson.
ITV4|1464041100|FYI Daily|23/05/2016||0|0|News Magazine,Current Affairs|
ITV4|1464041400|Heartbreak Ridge||1986|0|0|Adventure,War|A hellraising US marine sergeant is assigned to whip a squad of raw recruits into shape for the invasion of Grenada in 1983 - but his old-fashioned methods meet with disapproval from superior officers. Action adventure, directed by and starring Clint Eastwood. With Marsha Mason, Everett McGill, Moses Gunn and Bo Svenson.
ITV4|1464046800|Premiership Rugby Union|2015/16 Semi-Finals||0|0|Rugby Union - Domestic|Mark Durden-Smith and David Flatman present highlights of the semi-finals, which were Saracens v Leicester Tigers at Allianz Park and Exeter Chiefs v Wasps at Sandy Park.(n)
ITV4|1464050700|Motorsport UK|2016 Donington Park||0|0|Motor Sport|Action from Donington Park, featuring the MSA Formula Championship and the Ginetta GT4 Supercup. Commentary by Richard John Neil.(n)
ITV4|1464054300|ITV4 Nightscreen|||0|0|General Education,Science|Text-based information service.(n)
ITV4|1464055200|Teleshopping|||0|0|Advertisement,Shopping|Buying goods from the comfort of home.(n)
ITV4|1464066000|Hat-Trick Heroes|||0|0|General Sports|Short film featuring three-goal football heroes.(n)
ITV4|1464067200|Minder|You Gotta Have Friends||1|11|General Movie,Drama|Bearer bonds go missing from gangster Bobby Altman, and suspect Billy Gilpin appears at Arthur's house wanting to get out of town. Terry drives him to a hotel, but when Altman finds out he believes Arthur is involved and tries to establish the truth. George Baker and Roy Kinnear guest star.(n)
ITV4|1464071400|The Chase|24/05/2016||0|0|Quiz Show|Bradley Walsh presents as four contestants pit their wits against ruthless quiz genius the Chaser in the hope of winning a potential prize pot worth thousands of pounds. They work as a team and play strategically to answer general knowledge questions against the clock and race down the game board to the exit without being caught.(n)
ITV4|1464074700|MotoGP Highlights|2016 Italian Grand Prix||0|0|Motorcycling|The Italian Grand Prix. Action from the sixth round of the season, which was staged at the Mugello Circuit in Tuscany, Italy.(n)
ITV4|1464078600|Live French Open Tennis|2016 Day Three||0|0|Tennis|The third day of the Grand Slam tournament gets under way at Roland Garros, where more first-round matches are set to take place. Andy Murray began his campaign at last year's tournament with a straight-sets victory over `lucky loser' Facundo Arguello, while their were mixed fortunes for the two British ladies at the tournament, as Heather Watson defeated French wildcard entry Mathilde Johansson, but Johanna Konta lost to Denisa Allertova of the Czech Republic. Presented by John Inverdale, with analysis from Marion Bartoli, Jim Courier, Mark Petchey, Fabrice Santoro and Sam Smith, commentary by Nick Mullins and reports from Celina Hinchcliffe.(n)
ITV4|1464120000|The Chronicles of Riddick||2004|0|0|Adventure|Fugitive Riddick evades capture by bounty hunters and steals their spacecraft, only to run into an even bigger threat - fanatical cult members on a sinister mission to kill or convert anyone who crosses their path as they seek galactic domination. Sci-fi adventure sequel, with Vin Diesel reprising his role from Pitch Black alongside Judi Dench, Alexa Davalos and Thandie Newton.(n)
ITV4|1464123600|FYI Daily|24/05/2016 - 1||0|0|News Magazine,Current Affairs|
ITV4|1464123900|The Chronicles of Riddick||2004|0|0|Adventure|Fugitive Riddick evades capture by bounty hunters and steals their spacecraft, only to run into an even bigger threat - fanatical cult members on a sinister mission to kill or convert anyone who crosses their path as they seek galactic domination. Sci-fi adventure sequel, with Vin Diesel reprising his role from Pitch Black alongside Judi Dench, Alexa Davalos and Thandie Newton.(n)
ITV4|1464128400|30 Days of Night||2007|0|0|Horror|A horde of vampires finds the perfect hunting ground - a town in Alaska that remains sunless for a month. The local sheriff heads up a small band of townsfolk as they try to avoid the bloodthirsty invaders and survive until the sun rises once again. Horror, starring Josh Hartnett, Danny Huston and Melissa George.(n)
CITV|1463893200|The Aquabats! Super Show|Ladyfingers!||1|5|Cartoons,Puppets|The friends save a group of partying beachgoers from the threat of laser-blasting mummies.
CITV|1463894700|Pat & Stan|The Death of Norbert||1|10|Cartoons,Puppets|Pat and Stan decide to go to the seaside for the weekend with Stephanie, but at the last minute Stan realises he has forgotten Norbert, his stuffed animal.
CITV|1463895300|Dino Dan|There's a Compsognathus Under My Bed||1|5|General Children's,Youth|It is bedtime, but Dan is more interested in proving that there is a Compsognathus under his bed than going to sleep.
CITV|1463895900|Dino Dan|Art for Pterosaur's Sake||1|6|General Children's,Youth|Palaeontologist Dan Henderson and his friends make a kite inspired by the Quetzalcoatlus - but it remains to be seen whether it will fly.
CITV|1463896800|Signed Stories|Signed Stories: Share a Story: A Button||0|0|General Children's,Youth|A look behind the scenes of the Share a Story competition, meeting the competitors and the animators who turned their stories into short films.
CITV|1463897100|Sooty|The Rainy Day||2|15|General Children's,Youth|Heavy rain closes the park and leaks in the caravan roof, but expert plumbers Sooty and Sweep try to solve the problem.
CITV|1463897700|Super 4|A Colossal Challenge||1|9|Cartoons,Puppets|Animated comedy adventure series featuring a gang of heroes who protect the city of Technopolis and its King Kenric against evil elements.
CITV|1463898600|Nerds & Monsters|Hero Zeroes||1|16|Cartoons,Puppets|The children acquire superpowers after being bitten by a four-headed snake.
CITV|1463899500|The Tom & Jerry Show|Black Cat||1|46|General Children's,Youth|Madcap slapstick and mayhem as the celebrated cat and mouse plot against each other.
CITV|1463900400|Teen Titans Go|Let's Get Serious/Tamaranian Vacation||2|0|Cartoons,Puppets|The teenage superheroes fight to save the world while getting up to mischievous antics.
CITV|1463901900|Almost Naked Animals|Howie's Little Helper||1|52|General Children's,Youth|Chesley spends time with Howie for a school project, having decided to focus his attention on a hotel manager.
CITV|1463902800|Almost Naked Animals|Horn Swoggled||2|1|General Children's,Youth|Narwhal loses his horn, the source of his musical mojo, and switches jobs with Duck.
CITV|1463903700|Almost Naked Animals|The Night Shift||2|2|General Children's,Youth|Howie discovers there is a night shift at the Banana Cabana and that they have a lot more fun.
CITV|1463904600|Almost Naked Animals|The Green Banana||2|4|General Children's,Youth|Howie attempts to go green, but takes things too far.
CITV|1463905500|Almost Naked Animals|Trash in the Past||2|3|General Children's,Youth|Rubbish starts falling from the sky, prompting Howie and the gang to investigate.
CITV|1463906400|Almost Naked Animals|Howie's Pet Project||2|6|General Children's,Youth|Bunny challenges Howie to look after a pineapple for an entire afternoon.
CITV|1463907300|Almost Naked Animals|Dr Howie and Mr Howyena||2|5|General Children's,Youth|Howie creates a potion that turns him into an obnoxious party animal.
CITV|1463908200|Almost Naked Animals|Needle Day||2|8|General Children's,Youth|Children's entertainment.
CITV|1463909100|Almost Naked Animals|The Brother and Sister Games||2|9|General Children's,Youth|Howie makes a bet with Poodle that, if she can compete with him in The Brother and Sister Games, she can have half the hotel.
CITV|1463910000|Almost Naked Animals|Freebies Jeebies||2|10|General Children's,Youth|Howie sells coupons for the Banana Cabana, but Poodle doesn't like it as it's stealing her guests.
CITV|1463910900|Almost Naked Animals|Howie's Staycation||2|11|General Children's,Youth|Howie decides to take a staycation at the Banana Cabana by dressing up as a moose, but soon he meets a real version - who wants revenge on him.
CITV|1463911800|Almost Naked Animals|A Helping Paw||2|12|General Children's,Youth|Duck becomes Sloth's personal assistant when she only wants to spend time with Howie.
CITV|1463912700|Almost Naked Animals|Octo P.I.||2|13|General Children's,Youth|Octo discovers a real mystery while writing his novel.
CITV|1463913600|Almost Naked Animals|The Lost Stunt||2|14|General Children's,Youth|Howie tries to prove he is Dirk Danger's number one fan.
CITV|1463914500|City Shorts|Lights, Camera, Fire||1|4|Cartoons,Puppets|Children's game show.
CITV|1463914800|The Munch Box|||0|0|General Children's,Youth|Children's food challenge in which contestants battle it out to see who can come up with the most spectacular meal.
CITV|1463918400|House of Anubis|House of Heroes||3|40|General Children's,Youth|Eddie and KT try to unlock the portal and destroy Ammut once and for all. Alfie has a special gift for Willow.
CITV|1463919900|Oddbods|Hard and Heavy||1|35|General Children's,Youth|
CITV|1463920200|Fort Boyard Ultimate Challenge|Yellow Scorpions v Blue Sharks||4|1|Games and Quizzes|Adventure game show, in which teenage contestants from the UK and America compete in a series of quests around a fortress as they try to uncover hidden treasures. Presented by Laura Hamilton and Geno Segers.
CITV|1463922000|Fort Boyard Ultimate Challenge|Red Vipers v Silver Dragons||4|3|Games and Quizzes|The Red Vipers take on the Silver Dragons in the game show, in which teenage contestants compete in a series of quests around a fortress as they try to uncover hidden treasures. Presented by Laura Hamilton and Andy Akinwolere.
CITV|1463923500|City Shorts|Gold Run||0|0|Cartoons,Puppets|Children's game show.
CITV|1463923800|My Parents Are Aliens|Age Concerns||5|1|Comedy|Josh's voice breaks, making Brian and Sophie decide it's high time they started ageing too. Comedy, starring Danielle McCormack, Alex Kew and Charlotte Francis.
CITV|1463925600|Thunderbirds Are Go|Falling Skies||1|14|Cartoons,Puppets|Brains's latest invention - a self-constructing luxury space hotel - begins to malfunction, and International Rescue are called in to help.
CITV|1463927400|Grizzly Tales for Gruesome Kids|The New Nanny||1|1|General Children's,Youth|The cautionary story of two spoilt brats who meet their match in a nanny determined not to take any nonsense from them. Nigel Planer narrates.
CITV|1463928300|Grizzly Tales for Gruesome Kids|The Spaghetti Man||1|2|General Children's,Youth|Mirth and mayhem for younger viewers, based on the books by Jamie Rix and narrated by Nigel Planer.
CITV|1463929200|Horrid Henry|Horrid Henry and the Birthday Present||2|43|Cartoons,Puppets|Aunt Ruby takes Henry, Peter and Steve shopping for Mum's birthday present.
CITV|1463930100|Horrid Henry|Horrid Henry and the Zombie Hamster||2|44|Cartoons,Puppets|The mischievous boy's hamster Fang disappears and no-one knows if it is coming back.
CITV|1463931000|Horrid Henry|Horrid Henry Takes a Shortcut||2|40|Cartoons,Puppets|The friends discover that taking shortcuts will not always get you to your destination any quicker.
CITV|1463931900|Horrid Henry|Horrid Henry and the Antique Rogue Show||2|47|Cartoons,Puppets|The mischievous youngster and his friends discover that one person's rubbish is another's treasure.
CITV|1463932500|City Shorts|Lights, Camera, Fire||1|4|Cartoons,Puppets|Children's game show.
CITV|1463932800|Nerds & Monsters|Fab Rick||1|25|Cartoons,Puppets|An inflatable moose washes ashore, and Zarg destroys it.
CITV|1463934000|Nerds & Monsters|Inside the Box||1|26|Cartoons,Puppets|The children try to find out what is contained inside a strange crate.
CITV|1463934600|Almost Naked Animals|Howie Day||3|20|General Children's,Youth|Howie tries to complete enough good deeds to convince the mayor that he is worthy of his own special day.
CITV|1463935500|Almost Naked Animals|It's Duck's Party||3|22|General Children's,Youth|Narwhal has to keep Howie and the others from sneaking into Duck's very exclusive party.
CITV|1463936400|Deadtime Stories|Revenge of the Goblins||1|8|General Children's,Youth|Nina and Sammy release the goblins from under the earth - and now the repressed creatures are out for revenge.
CITV|1463937900|Signed Stories|Signed Stories: Share a Story: A Button||0|0|General Children's,Youth|A look behind the scenes of the Share a Story competition, meeting the competitors and the animators who turned their stories into short films.
CITV|1463938200|Looped|Baby Daddy||1|23|General Children's,Youth|Theo accidentally puts on anti-ageing cream and wakes to discover he is quickly ageing backwards.
CITV|1463939100|Looped|Wizard of Whacker Maze||1|24|General Children's,Youth|The school turns into a giant pinball game when Luc tries to defeat Kyle's high score.
CITV|1463940000|Horrid Henry|Horrid Henry's School Play||2|2|Cartoons,Puppets|The youngster has the chance to star in the school play, but has a good reason not to take the part.
CITV|1463940900|Horrid Henry|Horrid Henry and the Gross DVD||2|11|Cartoons,Puppets|Ralph lends Henry an unpleasant DVD, which the mischievous youngster cannot bring himself to watch.
CITV|1463941800|Thunderbirds Are Go|Falling Skies||1|14|Cartoons,Puppets|Brains's latest invention - a self-constructing luxury space hotel - begins to malfunction, and International Rescue are called in to help.
CITV|1463943600|Fort Boyard Ultimate Challenge|Yellow Scorpions v Blue Sharks||4|1|Games and Quizzes|Adventure game show, in which teenage contestants from the UK and America compete in a series of quests around a fortress as they try to uncover hidden treasures. Presented by Laura Hamilton and Geno Segers.
CITV|1463945400|Fort Boyard Ultimate Challenge|Red Vipers v Silver Dragons||4|3|Games and Quizzes|The Red Vipers take on the Silver Dragons in the game show, in which teenage contestants compete in a series of quests around a fortress as they try to uncover hidden treasures. Presented by Laura Hamilton and Andy Akinwolere.
CITV|1463946600|Oddbods|Critters and Cuisines||1|9|General Children's,Youth|The Oddbods have always had rather complicated relationships with animals, but their relationship with food is a lot simpler.
CITV|1463979600|Fleabag Monkeyface|Captain Maggotman||1|18|Cartoons,Puppets|Comic fans arrive for a convention, but the robotic Revoltoman goes out of control and kidnaps a famous inventor.
CITV|1463980200|Horrid Henry|Horrid Henry Says Goodbye||2|52|Cartoons,Puppets|The youngster has to move to another part of the country when his dad gets a new job, but decides to launch a counter campaign.
CITV|1463981100|Horrid Henry|Horrid Henry and the Gross Question||2|42|Cartoons,Puppets|The youngster searches for the answer to the `gross question', which lies in the most unexpected of places.
CITV|1463982000|Horrid Henry|Horrid Henry and the Birthday Present||2|43|Cartoons,Puppets|Aunt Ruby takes Henry, Peter and Steve shopping for Mum's birthday present.
CITV|1463982900|Matt Hatter Chronicles|Forest of Fears||3|9|General Children's,Youth|Matt, Roxie and Gomez battle two deadly foes - the Fire Phoenix and the bull-headed Minotaur - as Tenoroc tries to bend the inhabitants of the Enchanted Forest to his will.
CITV|1463984400|Matt Hatter Chronicles|Lightning Strikes Twice||3|10|General Children's,Youth|When a meteor storm splits Captain Lightning into two Captain Lightnings, Tenoroc pits the pair of livewires against each other to find some Multivisium ore for his masterplan.
CITV|1463986200|Thunderbirds Are Go|Designated Driver||1|22|Cartoons,Puppets|Alan's driving lessons with Parker take a much more urgent turn when burglars kidnap Lady Penelope and Aunt Sylvia. Action adventure, with the voices of Rasmus Hardiker, David Graham, Rosamund Pike and Sylvia Anderson.
CITV|1463987700|Almost Naked Animals|Life Was A Beach||0|0|General Children's,Youth|Children's animation featuring creatures who have shaved off their fur and wear only underclothes.
CITV|1463988600|Almost Naked Animals|Cabana Manana||1|51|General Children's,Youth|Howie trades away the beach, yard and pool in exchange for gifts for the others.
CITV|1463989500|Looped|Applecrab-dabra||1|11|General Children's,Youth|Animated adventures. Principal Applecrab's magic skills are put to the test when the boys cause a glitch and a real magician, Tommy Sparkles, shows up.
CITV|1463990400|Looped|Monday Circles||1|12|General Children's,Youth|Animated series following the adventures of two friends, Luc and Theo. Amy discovers the loop and spoils Luc and Theo's fun.
CITV|1463991000|Grizzly Tales for Gruesome Kids|Athlete's Foot||4|11|General Children's,Youth|A pair of ordinary-seeming running shoes hide a sinister secret dating from World War Two. Narrated by Nigel Planer.
CITV|1463991900|Grizzly Tales for Gruesome Kids|Grass Monkey||4|12|General Children's,Youth|Poor Spike falls in love with a girl who cares for her hair more than him. Narrated by Nigel Planer.
CITV|1463992800|Grizzly Tales for Gruesome Kids|The Top Hat||4|8|General Children's,Youth|A boy abuses the power of a magic hat, but is taught a lesson when the object swallows him and refuses to let him go.
CITV|1463993400|Sooty|It's a Dog's Life||2|19|General Children's,Youth|Sweep learns a valuable lesson in not taking his friends for granted as he realises there really is no place like home.
CITV|1463994300|Signed Stories|Signed Stories: Share a Story: The Donkey Tooth Fairy||0|0|General Children's,Youth|A look behind the scenes of the Share a Story competition, meeting the competitors and the animators who turned their stories into short films.
CITV|1463994600|Pat & Stan|Micro-Stan||1|23|Cartoons,Puppets|Stan the dog has a meeting with Professor Chi Chi.
CITV|1463995200|Pat & Stan|Bengal Hamster||1|24|Cartoons,Puppets|Stephanie and Pat offer Stan the dog a hamster to help calm him down.
CITV|1463995800|Dino Dan|Gasosaurus||1|10|General Children's,Youth|Dan Henderson and his friends learn that dino gas might have helped cause the extinction of the dinosaurs and cannot wait to share that information with the class.
CITV|1463996700|Dino Dan|He Shoots, He Roars||1|11|General Children's,Youth|Jim the reptile and his puppet Denny the dromaeosaurus help Dan figure out whether dinosaurs were warm-blooded.
CITV|1463997300|City Shorts|Adventures in the Air||1|2|Cartoons,Puppets|Children's game show.
CITV|1463997600|Super 4|Haunted Castle||1|12|Cartoons,Puppets|A ghost appears in the castle during Dr X's first visit to King Kenric, so Alex and his friends must do everything they can to get rid of it.
CITV|1463998500|Oddbods|A Day in the Life of Slick||1|5|General Children's,Youth|Slick is very tech-savvy and really cool, and he is mostly seen moving to a beat that is only in his head. Animated series.
CITV|1463998800|Oddbods|A Day in the Life of Bubbles||1|7|General Children's,Youth|Bubbles is the hungry yellow Oddbod, always optimistic and with a strange appetite for everything that moves. Animated series.
CITV|1463999400|Nerds & Monsters|It's Not Good to Be King||2|5|Cartoons,Puppets|Animated comedy about a group of children exiled on an uncharted island, where they have to be smart if they are to survive relentless attacks by a tribe of hideous monsters.
CITV|1464000300|Horrid Henry|Horrid Henry Says Goodbye||2|52|Cartoons,Puppets|The youngster has to move to another part of the country when his dad gets a new job, but decides to launch a counter campaign.
CITV|1464001200|Horrid Henry|Horrid Henry and the Gross Question||2|42|Cartoons,Puppets|The youngster searches for the answer to the `gross question', which lies in the most unexpected of places.
CITV|1464002100|Horrid Henry|Horrid Henry's Movie Moments||4|29|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.
CITV|1464003000|Horrid Henry|Hashtag Henry||4|25|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.
CITV|1464003900|Horrid Henry|Horrid Henry Goes on Strike||4|26|Cartoons,Puppets|Cartoon about a mischievous youngster. When Henry decides to go on strike, no-one is prepared for what happens.
CITV|1464004800|Horrid Henry|Moody Margaret for President||4|17|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.
CITV|1464005700|Fort Boyard Ultimate Challenge|Green Dragons vs White Falcons||0|0|Games and Quizzes|Adventure game show, in which teenage contestants from the UK and America compete in a series of quests around a fortress as they try to uncover hidden treasures.
CITV|1464007500|Fort Boyard Ultimate Challenge|Final Tournament||0|0|Games and Quizzes|Adventure game show, in which teenage contestants from the UK and America compete in a series of quests around a fortress as they try to uncover hidden treasures.
CITV|1464009000|Oddbods|Hard and Heavy||1|35|General Children's,Youth|
CITV|1464009300|Looped|The Replacements||1|13|General Children's,Youth|Animated series following the adventures of two friends. Luc and Theo vow to dethrone Sarah by taking over from Kelli and Kelly as her henchmen.
CITV|1464010200|Looped|Luc at Me||1|14|General Children's,Youth|Animated series following the adventures of two friends, Luc and Theo. In this edition, Luc enters a stunt contest.
CITV|1464011100|Almost Naked Animals|Horn Swoggled||2|1|General Children's,Youth|Narwhal loses his horn, the source of his musical mojo, and switches jobs with Duck.
CITV|1464012000|Almost Naked Animals|The Night Shift||2|2|General Children's,Youth|Howie discovers there is a night shift at the Banana Cabana and that they have a lot more fun.
CITV|1464012600|Dino Dan|A Winter Tail||1|12|General Children's,Youth|Trek wants to see some snow, but Dan Henderson is more concerned with seeing a euoplocephalus use its powerful tail.
CITV|1464013500|Dino Dan|Pterosaur in the House||1|13|General Children's,Youth|Ten-year-old Trek becomes obsessed with dinosaurs - and finds them everywhere.
CITV|1464014400|Super 4|Tower Trouble||1|13|Cartoons,Puppets|The heroes visit the castle and discover that Princess Leonora has been kidnapped, and set out to free her and also Ruby, who gets locked in the castle's keep.
CITV|1464015600|Nerds & Monsters|Tickle Stick||2|11|Cartoons,Puppets|When Becky is accidentally zapped by an electric sea creature, her braces light up and the Monsters begin using her for their various electrical needs.
CITV|1464016500|Nerds & Monsters|The Clown of Darkness||2|12|Cartoons,Puppets|Dudley discovers that comedy is an ideal way to distract the Monsters from eating the nerds, but takes his clowning a step too far.
CITV|1464017100|City Shorts|Adventures in the Air||1|2|Cartoons,Puppets|Children's game show.
CITV|1464017400|Mr Bean: The Animated Series|Super Trolley||1|29|Cartoons,Puppets|Faced with a long shopping list from his formidable landlady, the hapless half-wit builds a giant motorised trolley from a petrol mower and pram wheels, hoping to get the job done in double-quick time.
CITV|1464018300|Mr Bean: The Animated Series|Magpie||1|30|Cartoons,Puppets|The police suspect Bean of stealing his landlady's jewellery - but the real culprit is a magpie he's been nursing back to health.
CITV|1464019200|Looped|The Gifted Class||1|17|General Children's,Youth|Animated series. Luc and Theo discover a secret group for gifted kids and Theo is determined to join them.
CITV|1464020100|Looped|Sooper Loopers||1|18|General Children's,Youth|Animated adventures. The boys become superheroes.
CITV|1464021000|Adventure Time|Food Chain||6|7|General Children's,Youth|Finn goes on adventures with Jake the dog.
CITV|1464021900|Adventure Time|James II||6|3|General Children's,Youth|Finn goes on adventures with Jake the dog.
CITV|1464022800|Thunderbirds Are Go|Designated Driver||1|22|Cartoons,Puppets|Alan's driving lessons with Parker take a much more urgent turn when burglars kidnap Lady Penelope and Aunt Sylvia. Action adventure, with the voices of Rasmus Hardiker, David Graham, Rosamund Pike and Sylvia Anderson.
CITV|1464024300|Almost Naked Animals|Cabana Manana||1|51|General Children's,Youth|Howie trades away the beach, yard and pool in exchange for gifts for the others.
CITV|1464025200|Almost Naked Animals|Howie's Little Helper||1|52|General Children's,Youth|Chesley spends time with Howie for a school project, having decided to focus his attention on a hotel manager.
CITV|1464026100|Horrid Henry|Horrid Henry's Movie Moments||4|29|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.
CITV|1464027000|Horrid Henry|Hashtag Henry||4|25|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.
CITV|1464027900|Horrid Henry|Horrid Henry Goes on Strike||4|26|Cartoons,Puppets|Cartoon about a mischievous youngster. When Henry decides to go on strike, no-one is prepared for what happens.
CITV|1464028800|Horrid Henry|Moody Margaret for President||4|17|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.
CITV|1464029700|Oddbods|The Good, The Bad and the Insufferably Annoying||1|10|General Children's,Youth|Jeff snaps a winning photograph, Fuse races like a pro, and Pogo is the obnoxious prankster he normally is.
CITV|1464030000|Oddbods|Transportation Troubles||1|11|General Children's,Youth|The Oddbods share the many problems they encounter while using public transport.
CITV|1464030600|Nerds & Monsters|Monster Island: The Game||2|6|Cartoons,Puppets|Animated comedy about a group of children exiled on an uncharted island, where they have to be smart if they are to survive relentless attacks by a tribe of hideous monsters.
CITV|1464031500|Mr Bean: The Animated Series|Super Trolley||1|29|Cartoons,Puppets|Faced with a long shopping list from his formidable landlady, the hapless half-wit builds a giant motorised trolley from a petrol mower and pram wheels, hoping to get the job done in double-quick time.
CITV|1464032400|Mr Bean: The Animated Series|Magpie||1|30|Cartoons,Puppets|The police suspect Bean of stealing his landlady's jewellery - but the real culprit is a magpie he's been nursing back to health.
CITV|1464033300|Signed Stories|Signed Stories: Share a Story: When Some Aliens Came to My School||0|0|General Children's,Youth|Enchanting tales are conjured up from the magical Story Tree.(n)
CITV|1464066000|Fleabag Monkeyface|Raining Cats and Bogs||1|19|Cartoons,Puppets|A series of bizarre weather events have hit the city as it has been raining snails, snowing dandruff and gusting gales of boiled cabbage.(n)
CITV|1464066600|Horrid Henry|Horrid Henry and the Zombie Hamster||2|44|Cartoons,Puppets|The mischievous boy's hamster Fang disappears and no-one knows if it is coming back.(n)
CITV|1464067500|Horrid Henry|Horrid Henry Takes a Shortcut||2|40|Cartoons,Puppets|The friends discover that taking shortcuts will not always get you to your destination any quicker.(n)
CITV|1464068400|Horrid Henry|Horrid Henry and the Antique Rogue Show||2|47|Cartoons,Puppets|The mischievous youngster and his friends discover that one person's rubbish is another's treasure.(n)
CITV|1464069300|Matt Hatter Chronicles|The Tiger's Eye||3|11|General Children's,Youth|Tenor discovers that Roxie's staff can access great power at a place in the Enchanted Forest called the Neverglade, known only to Trackers.(n)
CITV|1464070800|Matt Hatter Chronicles|Shrinking Gas||3|12|General Children's,Youth|Tenor sends his latest super villain Gangster Bug into the critical airways that run under the Enchanted Forest.(n)
CITV|1464072600|Thunderbirds Are Go|Chain of Command||1|23|Cartoons,Puppets|Colonel Janus imposes a strict set of restrictions on the Thunderbirds after a series of mishaps nearly ends in disaster during a joint operation.(n)
CITV|1464074100|Almost Naked Animals|Horn Swoggled||2|1|General Children's,Youth|Narwhal loses his horn, the source of his musical mojo, and switches jobs with Duck.(n)
CITV|1464075000|Almost Naked Animals|The Night Shift||2|2|General Children's,Youth|Howie discovers there is a night shift at the Banana Cabana and that they have a lot more fun.(n)
CITV|1464075900|Looped|The Replacements||1|13|General Children's,Youth|Animated series following the adventures of two friends. Luc and Theo vow to dethrone Sarah by taking over from Kelli and Kelly as her henchmen.(n)
CITV|1464076800|Looped|Luc at Me||1|14|General Children's,Youth|Animated series following the adventures of two friends, Luc and Theo. In this edition, Luc enters a stunt contest.(n)
CITV|1464077400|Grizzly Tales for Gruesome Kids|Bugaboo Bear||0|0|General Children's,Youth|Mirth and mayhem for younger viewers, based on the books by Jamie Rix and narrated by Nigel Planer.(n)
CITV|1464078300|Grizzly Tales for Gruesome Kids|The Butcher Boy||5|2|General Children's,Youth|A boy's jealousy prompts him to steal the butcher's son's bike, but his actions lead to him finding out what it's like to be part of the meat industry.(n)
CITV|1464079200|Grizzly Tales for Gruesome Kids|The Fruit Bat||5|3|General Children's,Youth|A fussy girl learns about healthy eating the hard way when she is turned into a fruit bat.(n)
CITV|1464079800|Sooty|Record Breakers||2|20|General Children's,Youth|The puppet pals attempt to break world records for judge Boris McSquirter. Sooty tries to build a giant tower, while Sweep aims to become the world's tallest dog.(n)
CITV|1464080700|Signed Stories|Signed Stories: Share a Story: When Some Aliens Came to My School||0|0|General Children's,Youth|Enchanting tales are conjured up from the magical Story Tree.(n)
CITV|1464081000|Pat & Stan|In Search of Lost Treasure||1|25|Cartoons,Puppets|Aunt Martha comes across a strange map in an antique store which may lead to secret lost treasures.(n)
CITV|1464081600|Pat & Stan|Nasalation||1|26|Cartoons,Puppets|Stan grabs Pat's new perfume spray when it is delivered by the postman, but advertising claims that everyone will fall in love with whoever wears the scent soon prove to be untrue.(n)
CITV|1464082200|Dino Dan|A Winter Tail||1|12|General Children's,Youth|Trek wants to see some snow, but Dan Henderson is more concerned with seeing a euoplocephalus use its powerful tail.(n)
CITV|1464083100|Dino Dan|Pterosaur in the House||1|13|General Children's,Youth|Ten-year-old Trek becomes obsessed with dinosaurs - and finds them everywhere.(n)
CITV|1464083700|City Shorts|Fishing for Trouble||1|3|Cartoons,Puppets|Children's game show.(n)
CITV|1464084000|Super 4|Tower Trouble||1|13|Cartoons,Puppets|The heroes visit the castle and discover that Princess Leonora has been kidnapped, and set out to free her and also Ruby, who gets locked in the castle's keep.(n)
CITV|1464084900|Oddbods|A Day in the Life of Zee||1|8|General Children's,Youth|
CITV|1464085200|Oddbods|Critters and Cuisines||1|9|General Children's,Youth|The Oddbods have always had rather complicated relationships with animals, but their relationship with food is a lot simpler.(n)
CITV|1464085800|Nerds & Monsters|Monster Island: The Game||2|6|Cartoons,Puppets|Animated comedy about a group of children exiled on an uncharted island, where they have to be smart if they are to survive relentless attacks by a tribe of hideous monsters.(n)
CITV|1464086700|Horrid Henry|Horrid Henry and the Zombie Hamster||2|44|Cartoons,Puppets|The mischievous boy's hamster Fang disappears and no-one knows if it is coming back.(n)
CITV|1464087600|Horrid Henry|Horrid Henry Takes a Shortcut||2|40|Cartoons,Puppets|The friends discover that taking shortcuts will not always get you to your destination any quicker.(n)
CITV|1464088500|Horrid Henry|Horrid Henry and the Catastrophic Cushion||4|28|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464089400|Horrid Henry|Horrid Henry's Birthday Bonanza||4|33|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464090300|Horrid Henry|Horrid Henry Helps Out||4|31|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464091200|Horrid Henry|Horrid Henry's Vile Vacation||4|30|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464092100|The Aquabats! Super Show|ManAnt||1|1|Cartoons,Puppets|Crash is captured by the maniacal ManAnt, who plans to cipher his growth power to create an army of giant ants.(n)
CITV|1464093900|The Aquabats! Super Show|Mysterious Egg||1|2|Cartoons,Puppets|The Aquabats find a large egg in the forest and decide to incubate it, unaware a mutant monster bird is about to hatch.(n)
CITV|1464095400|Oddbods|More Than Enough||1|36|General Children's,Youth|The Oddbods have personalities as distinct as their furry suits and no two are alike. Animated series.(n)
CITV|1464095700|Looped|Loop it Forward||1|15|General Children's,Youth|Animated adventures of two friends, Luc and Theo. The boys decide to share their loop luck with an unlucky boy at school.(n)
CITV|1464096600|Looped|Chick Magnet||1|16|General Children's,Youth|Animated adventures of two friends, Luc and Theo. Theo sets out to impress Gwyn with a loopy science experiment.(n)
CITV|1464097500|Almost Naked Animals|The Green Banana||2|4|General Children's,Youth|Howie attempts to go green, but takes things too far.(n)
CITV|1464098400|Almost Naked Animals|Trash in the Past||2|3|General Children's,Youth|Rubbish starts falling from the sky, prompting Howie and the gang to investigate.(n)
CITV|1464099000|Dino Dan|Model Dino||1|14|General Children's,Youth|Ten-year-old Trek becomes obsessed with dinosaurs - and finds them everywhere.(n)
CITV|1464099900|Dino Dan|Copy Dino||1|15|General Children's,Youth|Ten-year-old Trek becomes obsessed with dinosaurs - and finds them everywhere.(n)
CITV|1464100800|Super 4|Fog Over Kingsland||1|14|Cartoons,Puppets|Animated comedy adventure series featuring a gang of heroes who protect the city of Technopolis and its King Kenric against evil elements.(n)
CITV|1464102000|Nerds & Monsters|Monstarrrghs!||2|13|Cartoons,Puppets|Irwin is excited because it is Talk Like a Pirate Day, but when he goes overboard and begins to annoy the other Nerds, he discovers he cannot stop.(n)
CITV|1464102900|Nerds & Monsters|The Sky's the Limit||2|14|Cartoons,Puppets|Becky tries to prove to Dudley that she does not need his help when it comes to mechanical know-how. Meanwhile, Zarg has shrinking head disease.(n)
CITV|1464103500|City Shorts|Fishing for Trouble||1|3|Cartoons,Puppets|Children's game show.(n)
CITV|1464103800|Mr Bean: The Animated Series|Cat Sitting||1|31|Cartoons,Puppets|The fur flies when Scrapper is left in Mr Bean's care - and it's not the creepy cat who needs looking after in the end. With the voice of Rowan Atkinson.(n)
CITV|1464104700|Mr Bean: The Animated Series|The Bottle||1|32|Cartoons,Puppets|A milkman accidentally walks off with a maritime curio belonging to Bean - who indignantly follows him to the bottling plant at the local dairy, determined to retrieve it.(n)
CITV|1464105600|Almost Naked Animals|Trash in the Past||2|3|General Children's,Youth|Rubbish starts falling from the sky, prompting Howie and the gang to investigate.(n)
CITV|1464106500|Almost Naked Animals|Howie's Pet Project||2|6|General Children's,Youth|Bunny challenges Howie to look after a pineapple for an entire afternoon.(n)
CITV|1464107400|Adventure Time|The Red Throne||5|47|General Children's,Youth|Finn goes on adventures with Jake the dog.(n)
CITV|1464108300|Adventure Time|Betty||5|48|General Children's,Youth|Finn goes on adventures with Jake the dog.(n)
CITV|1464109200|Thunderbirds Are Go|Chain of Command||1|23|Cartoons,Puppets|Colonel Janus imposes a strict set of restrictions on the Thunderbirds after a series of mishaps nearly ends in disaster during a joint operation.(n)
CITV|1464110700|Almost Naked Animals|Horn Swoggled||2|1|General Children's,Youth|Narwhal loses his horn, the source of his musical mojo, and switches jobs with Duck.(n)
CITV|1464111600|Almost Naked Animals|The Night Shift||2|2|General Children's,Youth|Howie discovers there is a night shift at the Banana Cabana and that they have a lot more fun.(n)
CITV|1464112500|Horrid Henry|Horrid Henry and the Catastrophic Cushion||4|28|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464113400|Horrid Henry|Horrid Henry's Birthday Bonanza||4|33|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464114300|Horrid Henry|Horrid Henry Helps Out||4|31|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464115200|Horrid Henry|Horrid Henry's Vile Vacation||4|30|Cartoons,Puppets|Cartoon about a mischievous youngster who delights in playing pranks, being rotten to his relatives and generally getting up to no good.(n)
CITV|1464116100|Oddbods|Exercise Overload||1|12|General Children's,Youth|
CITV|1464116400|Oddbods|In For a Rocky Ride||1|13|General Children's,Youth|
CITV|1464117000|Nerds & Monsters|Nerd Fu||2|7|Cartoons,Puppets|Animated comedy about a group of children exiled on an uncharted island, where they have to be smart if they are to survive relentless attacks by a tribe of hideous monsters.(n)
CITV|1464117900|Mr Bean: The Animated Series|Cat Sitting||1|31|Cartoons,Puppets|The fur flies when Scrapper is left in Mr Bean's care - and it's not the creepy cat who needs looking after in the end. With the voice of Rowan Atkinson.(n)
CITV|1464118800|Mr Bean: The Animated Series|The Bottle||1|32|Cartoons,Puppets|A milkman accidentally walks off with a maritime curio belonging to Bean - who indignantly follows him to the bottling plant at the local dairy, determined to retrieve it.(n)
Channel 5|1463871600|SuperCasino|||0|0|Game Show,Quiz|Viewers get the chance to take part in live interactive gaming, with an entertaining mix of roulette-wheel spins and lively chat from the presenting team. Featuring a variety of prizes and promotions.
Channel 5|1463883000|Spike Fight Night|BAMMA 25: Champion vs Champion||0|0|Boxing|Action from the event staged at Barclaycard Arena in Birmingham, where three title bouts were set to take place, including Shay Walsh v Tom DuQuesnoy for the Bantamweight belt.
Channel 5|1463889300|Divine Designs|Temples of Suburbia||2|15|General Arts,Culture|Dr Paul Binski, Professor of the History of Medieval Art at Cambridge University, examines religious art, viewing spectacular Hindu and Jain works in Leicester and north London.
Channel 5|1463890800|House Doctor|Spennymoor||6|4|Property|Property guru Ann Maurice applies her home improvement remedies to a house in Spennymoor, Co Durham, for the purpose of finding an eager buyer as soon as possible.
Channel 5|1463892300|Angels of Jarm|Fatima's Mum||1|14|General Children's,Youth|Wendy is scared of Fatima's mum because of her clothes.
Channel 5|1463892600|Angels of Jarm|Don't Touch!||1|15|General Children's,Youth|The children are warned not to touch anything in the kitchen, but when they start baking cakes Angel Rafe has to come down and look after them.
Channel 5|1463893200|Peppa Pig|The Cycle Ride||2|33|Cartoons,Puppets|The family spends the day riding bikes, and participate in a downhill race.
Channel 5|1463893500|Bananas in Pyjamas|A Bunch of Bananas||2|44|Cartoons,Puppets|The duo are impressed with Charlie's latest invention - a super ball that never stops bouncing, but when they accidentally let it out of the workshop, they struggle to catch it. Animation, featuring the voices of Richard McCourt and Dominic Wood.
Channel 5|1463894100|Angelina Ballerina|Angelina's Rock Band||3|15|Cartoons,Puppets|The youngster's friends rehearse in a band for a school project and invite her to join in as the tambourine player.
Channel 5|1463895000|Bob the Builder|Out of the Woods||1|31|Cartoons,Puppets|Bob and the team work at Fixham campsite, where Leo alarms the machines with his spooky stories and Dizzy takes care of an injured creature.
Channel 5|1463895900|Tickety Toc|Fix-It Time||2|8|Cartoons,Puppets|McCoggins leaves the twins alone in his workshop, so Tommy decides to try to mend a broken truck, but forgets to put back an important red button.
Channel 5|1463896500|Zack and Quack|Pop-Up Speedway||1|6|Cartoons,Puppets|The gang builds a pop-up race car, and Zack wants to prove it can be a winner on the track.
Channel 5|1463897100|Pets|Kittens||1|9|General Children's,Youth|Two sisters make toy spiders for their kittens to play with, but have a hard time tempting their pets out from under the sofa.
Channel 5|1463897400|Noddy in Toyland|Tessie and the Fairy Cakes||1|40|General Children's,Youth|Tessie adds fairy powder to her cakes in an effort to gain an unfair advantage over Mr Wobbly Man in a baking contest.
Channel 5|1463898300|Paw Patrol|Pups and the Mischievous Kittens||2|18|Cartoons,Puppets|To win the Spotless Town award, the Paw Patrol pups must save Adventure Bay from Mayor Humdinger's kitten catastrophe crew.
Channel 5|1463899200|Little Princess|I Want My Robin||3|33|Cartoons,Puppets|The youngster goes bird-watching, but the wild creatures are difficult to see as they keep flying off.
Channel 5|1463899800|Pip Ahoy|The New Harbour Pilot||1|34|Cartoons,Puppets|Salty Cove needs a new harbour pilot, and Mr Morris would love the job, but thinks he might not be fit enough. Pip, Alba and friends decide to put him through his paces.
Channel 5|1463900700|Blaze and the Monster Machines|Cattle Drive||1|15|General Children's,Youth|Blaze and Starla find a herd of cows wandering in the desert, and set out to bring them back to Starla's barn.
Channel 5|1463902200|Ben and Holly's Little Kingdom|Gaston to the Rescue||2|15|General Children's,Youth|The elves and fairies encounter a speaking door and a dwarf mine while on the lookout for Gaston.
Channel 5|1463903400|Wanda and the Alien|Hiccups||1|35|General Children's,Youth|Daddy Rabbit makes some fizzy carrot juice that gives everyone a bad case of the hiccups, including the squirrels, so Wanda and Alien go in search of a cure.
Channel 5|1463904000|Toby's Travelling Circus|Plunger Fun||1|27|General Arts,Culture|Dolores takes a plunger Clara and Freddo have incorporated into their routine to unblock a sink in her caravan, but when she gets locked in, the gang races to return the tool to the duo in time for the show.
Channel 5|1463904900|Jelly Jamm|Apprentice Bello||1|21|General Children's,Youth|Apprentice Bello is put in charge of operating the Music Factory.
Channel 5|1463905800|LazyTown|Who's Who?||3|5|General Children's,Youth|Robbie Rotten dislikes Stephanie teaching everyone how to dance, and creates a robot clone of her that says discouraging things to the LazyTowners. The real Stephanie has to be discovered through a dance-off.
Channel 5|1463907300|Teenage Mutant Ninja Turtles|The Noxious Avenger||3|15|Animated Movie,Drama|A new mutant called Muckman starts gain notoriety as New York City's new `Monster Hero'.
Channel 5|1463909400|Now That's Funny|||1|3|Family|Amusing Internet-sourced videos, including pleasure seekers getting more than they bargained for at an amusement park and people who have turned fooling about at work into an art form. Plus, kung fu bears, screaming samurais and clumsy creatures.
Channel 5|1463912700|Cloudy with a Chance of Meatballs 2||2013|0|0|Animated Movie,Drama|A scientist believes he has saved the world from his invention, a machine that accidentally turned water into food. However, he learns the device is still active and has created a race of food/animal hybrids that he must stop from running wild across the world. Animated comedy sequel, with the voices of Bill Hader, Anna Faris and James Caan.
Channel 5|1463919000|Most Shocking Talent Show Moments|||0|0|Documentary|Countdown of 50 of the most memorable moments from TV talent shows, including Rylan's outrageous antics on The X Factor in 2012 and life-changing first appearances on Britain's Got Talent by Susan Boyle and Paul Potts. Featuring contributions by Anton Du Beke, Craig Revel Horwood, Ann Widdecombe, Matthew Kelly, Pete Waterman, Nicki Chapman and Eddie `the Eagle' Edwards.
Channel 5|1463929500|Pudsey the Dog: The Movie||2014|0|0|Comedy|Premiere. A stray dog who has always looked out for number one learns the benefits of having a family when he is adopted by a single mother and her three children in a sleepy seaside village. He realises his new owners' landlord is up to no good and tries to foil his evil plans. Family comedy, starring Jessica Hynes and John Sessions, with the voice of David Walliams.
Channel 5|1463936100|The Yorkshire Vet|||1|1|General Arts,Culture|Documentary about Yorkshire vet Julian Norton, his business partner Peter Wright and their team as they administer modern-day medical and surgical aid to creatures great and small. In the first episode, Julian treats a much-loved cat with a swollen eye, for which surgery might be the only option. He also steps in to find out what is wrong with Copper, Head Nurse Sarah's beloved dog.
Channel 5|1463939700|5 News Weekend|22/05/2016||0|0|News|Round-up of the day's headlines from around the world.
Channel 5|1463940000|Cricket on 5|England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. Highlights from the fourth day of the First Test in a three-match series, which takes place at Headingley. Presented by Mark Nicholas, who also commentates alongside Michael Vaughan, Geoffrey Boycott, and Simon Hughes.
Channel 5|1463943600|Secrets of Egypt|Secrets of the Valley of the Kings: Valley of the Kings||0|0|Documentary|An exploration of the Valley of the Kings, the royal necropolis of the pharaohs and the world's most famous royal burial ground. Egyptologists investigate what drove Egypt's greatest pharaohs to seek out this secluded valley to hide their remains, how ancient craftsmen managed to achieve such feats of engineering and keep pace with the ever-shifting designs, and why was the sacred site was finally abandoned. Narrated by Mark Halliley.
Channel 5|1463947200|Sabotage||2014|0|0|Police,Crime Drama|The members of an elite Drug Enforcement Administration team secretly keep the millions of dollars they find during the raid. When they are killed off one by one, the leader becomes convinced one of his men is getting rid of the others to keep all the money, and sets out to expose the murderer. Action thriller, starring Arnold Schwarzenegger and Sam Worthington.
Channel 5|1463954700|Under Siege||1992|0|0|Adventure|Terrorists infiltrate a US battleship in a carefully orchestrated move to steal its arsenal of nuclear weapons, unaware the ship's resourceful cook - a veteran US Navy Seal - and a scantily clad stripper are about to foil their plans. Action adventure, starring Steven Seagal, Erika Eleniak, Gary Busey and Tommy Lee Jones. Edited for broadcast.
Channel 5|1463961300|SuperCasino|||0|0|Game Show,Quiz|Viewers get the chance to take part in live interactive gaming, with an entertaining mix of roulette-wheel spins and lively chat from the presenting team. Featuring a variety of prizes and promotions.
Channel 5|1463969400|Police Interceptors|||10|10|Factual Crime|Paul Faulkner has a close shave with a stolen vehicle, Kev Salter takes part in a stake-out, Liam has a front-row seat in a pirouetting pursuit and Spike unearths a bumper crop of cannabis.
Channel 5|1463972400|Now That's Funny|||1|3|Family|Amusing Internet-sourced videos, including pleasure seekers getting more than they bargained for at an amusement park and people who have turned fooling about at work into an art form. Plus, kung fu bears, screaming samurais and clumsy creatures.
Channel 5|1463975400|Nick's Quest|Anaconda||1|1|Nature,Animals|Naturalist Nick Baker searches for the world's most dangerous animals. He begins with a trip to the remote Llanos region of Venezuela in the hope of encountering the anaconda, one of nature's largest snakes.
Channel 5|1463976900|Nick's Quest|Great White Shark||1|2|Nature,Animals|Nick Baker examines the habits of the great white shark, which can grow to 20ft in length. From the safety of an underwater cage, he has an encounter with one of the creatures off the Western Cape of South Africa. He also swims with fur seals and penguins.
Channel 5|1463978700|Angels of Jarm|Singing Angel||1|16|General Children's,Youth|The children worry about singing in class - until Angel Ellie arrives.
Channel 5|1463979000|Angels of Jarm|Symbols||1|17|General Children's,Youth|The children laugh at Aaron when he draws a star with six points.
Channel 5|1463979600|The WotWots|Topsy Turvy Wotty||1|20|Cartoons,Puppets|The aliens learn about creatures that hang upside down.
Channel 5|1463980200|Chloe's Closet|Turtle Fishing||2|21|General Children's,Youth|Chloe goes fishing and has to help a turtle that has lost its babies.
Channel 5|1463980800|Lily's Driftwood Bay|Message in a Bottle||1|23|Cartoons,Puppets|It's Gull's birthday and after Lily finds a message in a bottle on the beach, they have fun following a mysterious trail of clues around the bay.
Channel 5|1463981400|Fireman Sam|Open Day||6|25|Cartoons,Puppets|Pontypandy Fire Station is opened to the public and Norman is eager to try things out, crawling under safety tape and getting into the driving seat of a fire engine. However, his inquisitive nature and desire for excitement lead to danger when he climbs onto the roof to get closer to Tom and his helicopter.
Channel 5|1463982000|Wissper|Pig in a Puddle||1|15|Cartoons,Puppets|A mummy pig's piglets cannot cover themselves in mud because their waterhole has dried up.
Channel 5|1463982600|Peppa Pig|Fish Pond||4|48|Cartoons,Puppets|Daddy Pig takes Peppa and George to a fish pond that he used to visit when he was a piglet.
Channel 5|1463982900|Pip Ahoy|Bubble Trouble||1|35|Cartoons,Puppets|Alba and Pip volunteer to help Skipper wash up, and when Hopper is sent to get a fresh bottle of washing-up liquid, the whole of Salty Cove is mysteriously flooded with bubbles.
Channel 5|1463983800|Little Princess|I Want to Recycle||3|34|Cartoons,Puppets|The youngster realises the importance of not wasting things and tries to think of ways to recycle rubbish.
Channel 5|1463984400|Bob the Builder|Never Give Up||1|32|Cartoons,Puppets|While Bob and his team set to work on a new zipline, Leo makes mistakes and starts to question whether or not he is cut out to be a builder.
Channel 5|1463985300|Thomas & Friends|No Steam Without Coal||18|14|Cartoons,Puppets|Timothy warns Bill and Ben to use their coal sensibly when there is a shortage at the Clay Pits, but they choose not to listen to him and soon run out of fuel.
Channel 5|1463986200|Noddy: Toyland Detective|Noddy and the Case of the Sticky Putty||1|13|General Children's,Youth|Noddy realises that someone has put sticky putty on Clockwork Mouse's key, and comes up with a clever solution when he finds out who did it and why.
Channel 5|1463986800|Ben and Holly's Little Kingdom|Miss Cookie's Nature Trail||2|16|General Children's,Youth|Miss Cookie organises a nature trail for Lucy and her class, but it goes through the middle of the Little Kingdom.
Channel 5|1463987700|Peppa Pig|Dens||2|36|Cartoons,Puppets|Peppa announces only girls are allowed to play in her treehouse, so Grandpa Pig builds the boys their own den.
Channel 5|1463988300|Peppa Pig|Zoe Zebra the Postman's Daughter||2|28|Cartoons,Puppets|Zoe joins her postman dad Mr Zebra on his daily rounds.
Channel 5|1463988900|Paw Patrol|Pups Save a Friend||2|19|Cartoons,Puppets|When Marshall decides to take a break from the Paw Patrol, the pups jump into action to bring him back.
Channel 5|1463989800|Bananas in Pyjamas|The Banana Dance||2|45|Cartoons,Puppets|The duo want to make up a new dance to show everyone at the Cuddlestown dance party, but have to work on it quickly.
Channel 5|1463990400|Toot the Tiny Tugboat|Toot Needs Help||1|19|Cartoons,Puppets|Toot hopes to impress the admiral with his hard work - but he learns he cannot do everything by himself.
Channel 5|1463991300|The Wright Stuff|23/05/2016||0|0|Discussion,Debate|Journalist and broadcaster Matthew Wright is joined by a panel of guests and the studio audience to debate the issues of the day.
Channel 5|1463998500|GPs: Behind Closed Doors|||3|12|Medicine,Health|In this edition, the doctors at Balham Park Surgery must deal with several highly emotional patients. Dr Eleanor Beecraft's patient is furious that his ears are still blocked up with wax, despite him consistently missing hospital appointments to have them syringed. Meanwhile, a woman arrives for an appointment with Dr Shah, and is terrified that her stomach pains are a sign of ovarian cancer. Dr Heather Watson sees a patient who, instead of feeling ecstatic at being newly pregnant, is in mortal fear of another miscarriage.
Channel 5|1464001800|5 News Lunchtime|23/05/2016||0|0|News|Round-up of the day's headlines from around the world.
Channel 5|1464002100|Cowboy Builders & Bodge Jobs|Cowboy Builders||1|8|Property|Dan Lobb and Laura Hamilton travel to Newbury to meet Nicky, whose mother Jill took the opportunity to move into the house next door when it went up for sale. However, cracks began to appear after building work started, and Jill ended up with a toilet in her bedroom, facing the prospect of making trips to her daughter's to wash herself.
Channel 5|1464005700|Home and Away|||0|0|Soap,Melodrama|Sun-kissed Australian soap charting the latest comings and goings of the Summer Bay regulars.
Channel 5|1464007500|Neighbours|||0|0|Soap,Melodrama|Having learned the real identity of `Mitch', Sonya decides to confront Uncle Walter. Lauren doubts Brad's fidelity, while Piper unearths a new suspect for the Lassiter's blast.
Channel 5|1464009600|NCIS: New Orleans|Musician Heal Thyself||1|2|Detective,Thriller|A case becomes personal for Pride when a murder victim is identified as Petty Officer Calvin Parks, who the agent used to mentor when the young man was in a gang. LaSalle question members of two rival gangs, but a drive-by shooting linked to the killing leads to an accusation from a mayoral candidate that the NCIS team has stirred up violence, and the investigators begin to question whether the death has a political connection. Crime drama, starring Scott Bakula and Lucas Black.
Channel 5|1464012900|Killer Switch||2016|0|0|General Movie,Drama|A woman accidentally picks up the wrong suitcase from the airport baggage reclaim on her way to her daughter's graduation. Later, she receives a phone call from a man claiming he will harm her daughter if she fails to follow his instructions to return his suitcase. Thriller, starring Jamie Luner.
Channel 5|1464019200|5 News at 5|23/05/2016||0|0|News|Round-up of the day's headlines from around the world.
Channel 5|1464021000|Neighbours|||0|0|Soap,Melodrama|Having learned the real identity of `Mitch', Sonya decides to confront Uncle Walter. Lauren doubts Brad's fidelity, while Piper unearths a new suspect for the Lassiter's blast.
Channel 5|1464022800|Home and Away|||0|0|Soap,Melodrama|Sun-kissed Australian soap charting the latest comings and goings of the Summer Bay regulars.
Channel 5|1464024600|5 News Tonight|23/05/2016||0|0|General News,Current Affairs|A round-up of the evening's headlines, including coverage of the latest national and international stories.
Channel 5|1464026100|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Vote Leave campaign.
Channel 5|1464026400|Cricket on 5|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights from the fifth day of the First Test in a three-match series, which took place at Headingley. Presented by Mark Nicholas, who also commentates alongside Michael Vaughan, Geoffrey Boycott, and Simon Hughes.
Channel 5|1464030000|Police Interceptors|||10|11|Factual Crime|Chris and Andy pursue a drug dealer through the back streets of Shotton, Co Durham, Kev tracks down a man threatening drinkers with an axe, and Spike has a high-speed chase in the countryside. Finally, Richie learns that perseverance sometimes bring its own reward.
Channel 5|1464033600|Secrets of the Nazi Occult|||0|0|Documentary|Documentary examining a secret society that contained many members of the Nazi high command, including both Adolf Hitler and Heinrich Himmler, and which held meetings and conducted rituals at Wewelsburg Castle in Germany.
Channel 5|1464037200|Gotham|Gotham: Wrath of the Villains: Azrael||2|19|Detective,Thriller|Gordon questions Strange about Project Chimera and also serves a writ ordering an exhumation, which leads the professor to send the newly resurrected Galavan to deal with the detective. Meanwhile, Ed Nygma begins to understand how to manipulate his fellow inmates to get them on his side.
Channel 5|1464040800|Up Late with Rylan|||1|9|Talk Show|Rylan Clark-Neal hosts the chat show, featuring celebrity guests and music as well as games for the studio audience and the viewers at home.
Channel 5|1464043500|Nightmare Tenants, Slum Landlords|||2|11|Documentary|Claire and Simon seek eviction specialist Chris's help to evict a man claiming to be renting their old family home. Meanwhile, Hazma hopes to get his council flat back after he tried to help a neighbour's friend by letting them stay for a week, but ended up being shut out when they refused to leave. Plus, a man is almost £30k in debt and in danger of repossession after his tenants stopped paying the rent.
Channel 5|1464047100|Tattoo Disasters UK|||1|1|General Education,Science|People who regret their tattoos share the stories behind their body art and take steps to get them removed. A woman describes a desperate attempt to erase a former partner's name from her wrist, a man reveals how he woke from a wild night out with a slogan inked on his back and the most tattooed man in Britain reveals his latest addition. Plus, the aspiring model who now regrets getting a huge tattoo of a disgraced pop star on her stomach.(n)
Channel 5|1464048600|SuperCasino|||0|0|Game Show,Quiz|Viewers get the chance to take part in live interactive gaming, with an entertaining mix of roulette-wheel spins and lively chat from the presenting team. Featuring a variety of prizes and promotions.(n)
Channel 5|1464055800|Castle|Countdown||3|17|Detective,Thriller|Part two of two. Ryan and Esposito manage to track down Beckett and Castle to the freezer container and rescue them in the nick of time. Agent Fallon reinstates them after admitting they were on the right track in pursuit of the bomber threatening New York, and their investigation leads them to a woman who recognises the taxi driver as a man who served in the same regiment as her late brother Kevin.(n)
Channel 5|1464058800|Caught on Camera|Criminals: Caught on Camera||1|1|Factual Crime|Journalist Nick Wallis joins police forces across the nation to discover how CCTV and other technological advances are helping to bring criminals to justice. The first episode focuses on drunkenness and violence, with Nick going to Chester on a race day to find out how the local council and police are using cameras to deal with the 50,000 people descending on the city. In Rotherham, South Yorkshire, operators Martyn and Dave keep in radio contact with nightclub bouncers to prevent trouble at the weekend.(n)
Channel 5|1464061500|Wildlife SOS|||2|21|Nature,Animals|The work of volunteers treating sick, injured and orphaned animals at a wildlife sanctuary.(n)
Channel 5|1464063000|Great Artists|Leonardo||1|2|Fine Arts|Tim Marlow profiles scientist, engineer, inventor and painter Leonardo da Vinci, whose extraordinary artistic genius gave rise to masterpieces including the Mona Lisa, the Annunciation and the Last Supper. Breaking new ground in portraiture and historical imagery, this giant of the Italian Renaissance used his wide-ranging skills to make a unique contribution to the development of European art.(n)
Channel 5|1464064500|House Doctor|Headcorn||2|2|Property|Ann Maurice visits Headcorn to help a couple spruce up their tiny cottage in a bid to make it more attractive to prospective buyers, clearing out all their clutter, getting rid of a dingy carpet and using small furniture to create an illusion of space.(n)
Channel 5|1464066000|The WotWots|Go the Greens||1|21|Cartoons,Puppets|SpottyWot refuses to eat broccoli soup, so DottyWot shows him that greens are important.(n)
Channel 5|1464066600|Chloe's Closet|A Super Sticky Situation||2|22|General Children's,Youth|Chloe and her friends develop super powers and must use them to save a carnival from a destructive pair of giant lobsters.(n)
Channel 5|1464067200|Lily's Driftwood Bay|Stop! Watch||1|24|Cartoons,Puppets|Lily finds Salty's pocket watch, but has it snatched from her by the Clickety Clackety train.(n)
Channel 5|1464067800|Fireman Sam|Mike's Rocket||6|26|Cartoons,Puppets|Norman tries to produce a spectacle to rival Mike's rocket show by holding his own in Pontypandy.(n)
Channel 5|1464068400|Wissper|Thirsty Giraffe||1|16|Cartoons,Puppets|Gertie the giraffe needs help bending down to take a drink, so Wissper enlists the help of Peggy the penguin to raise the water level.(n)
Channel 5|1464069000|Peppa Pig|The Olden Days||4|51|Cartoons,Puppets|Mummy Pig shows Peppa and her friend Suzy Sheep some old photographs from when they were babies.(n)
Channel 5|1464069300|Pip Ahoy|The Alan Comet||1|36|Cartoons,Puppets|A comet is due to fly over Salty Cove and everyone wants to stay awake to see it. Hopper decides to have a nap during the day so he can stay up all night - but his rest is disturbed by Alan the Penguin.(n)
Channel 5|1464070200|Little Princess|Who Turned the Lights Off?||3|35|Cartoons,Puppets|The castle suffers a power cut just as the household is preparing for a birthday party.(n)
Channel 5|1464070800|Bob the Builder|Smallest Rocket||1|33|Cartoons,Puppets|Bob and the team are asked to build the launch pad for Mei Moon's rocket, but the launch is in danger of being cancelled when Lofty makes a mistake.(n)
Channel 5|1464071700|Thomas & Friends|Spencer's VIP||18|15|Cartoons,Puppets|Spencer brings a VIP back from the mainland, but arrives so late that the passenger refuses to travel with him. The other engines then compete to be chosen for the exciting task.(n)
Channel 5|1464072600|Noddy: Toyland Detective|Noddy and the Case of the Broken Crystal Memory Game'||1|1|General Children's,Youth|The DareDale Challenge obstacle race is about to start when it is discovered that the crystal memory game is broken. While Clockwork Mouse sets about mending it, Noddy and Revs try to find out who was responsible.(n)
Channel 5|1464073200|Ben and Holly's Little Kingdom|The New Wand||2|17|General Children's,Youth|Holly's wand catches a cold and she is given a WiseWand 3000 as a replacement.(n)
Channel 5|1464074100|Peppa Pig|The Cuckoo Clock||2|30|Cartoons,Puppets|Daddy Pig winds up the old cuckoo clock in Peppa and George's bedroom.(n)
Channel 5|1464074700|Peppa Pig|Ice Skating||2|34|Cartoons,Puppets|The friends go ice-skating, but keep falling over.(n)
Channel 5|1464075300|Paw Patrol|Pups Save a Stowaway||2|20|Cartoons,Puppets|When the pups find a stowaway on their trip to the icy tundra, they must rescue a runaway kitty on a runaway snowcat.(n)
Channel 5|1464076200|Bananas in Pyjamas|The Pen Pal||2|46|Cartoons,Puppets|Amy's pen pal is always telling her about all the amazing stuff he does, so the Bananas follow her and make a list of all the special things she does.(n)
Channel 5|1464076800|Toot the Tiny Tugboat|Flag Day||1|20|Cartoons,Puppets|Toot has not done much to prepare his contribution to Flag Day, and leaves everything until it is almost too late. He has to rush to finish, and learns the value of being organised.(n)
Channel 5|1464077700|The Wright Stuff|24/05/2016||0|0|Discussion,Debate|Matthew Wright and guests talk about the issues of the day, with viewers calling in to offer their opinions.(n)
Channel 5|1464084900|GPs: Behind Closed Doors|||3|13|Medicine,Health|Dr William Laird tries to help a patient suffering from chronic vertigo, twisting their head in an attempt to shift the debris inside the ear that is causing the problem. Meanwhile, Dr Shah gets busy with a tuning fork, pressing against a patient's skull to ascertain the severity of a man's debilitating tinnitus.(n)
Channel 5|1464088200|5 News Lunchtime|24/05/2016||0|0|News|Round-up of the day's headlines from around the world.(n)
Channel 5|1464088500|Cowboy Builders & Bodge Jobs|Cowboy Builders||1|9|Property|John Russell and Laura Hamilton travel to Mitcham, south London, to meet a couple who need help transforming their half-finished loft conversion into a bedroom. They started the project because they were desperate for their parents to have a place to stay so they could help raise their young daughter and newborn baby, but their builder failed to complete the job.(n)
Channel 5|1464092100|Home and Away|||0|0|Soap,Melodrama|Zac is forced to perform life-saving emergency surgery on Hunter, Skye teases VJ when she realises he has a crush on Billie, and Greg finds out Zac was in prison with his son Wayne.(n)
Channel 5|1464093900|Neighbours|||0|0|Soap,Melodrama|Brodie divulges a piece of detail regarding the Lassiter's blast that he should not know. Terese seeks distraction from her grief, while Lauren feels uneasy about Ned.(n)
Channel 5|1464095700|NCIS|We Build, We Fight||12|13|Detective,Thriller|Gibbs and his colleagues investigate when Eric Kutzler, the first openly gay Navy lieutenant tipped to receive the Medal of Honour, is murdered. While the agents initially suspect Kutzler's death was the result of a hate crime, the fact that his police officer husband waited 20 minutes to report the crime suggests he had something to hide. Meanwhile, the team throws a baby shower for Palmer as his wife's due date approaches. Starring Mark Harmon, Michael Weatherly and Pauley Perrette.(n)
Channel 5|1464099300|Seduced by Lies||2010|0|0|Thriller|A woman hopes to make a fresh start with a new relationship in defiance of her father's wishes, and turns her back on old friends when they are suspicious of her boyfriend. However, she gradually comes to realise that he has a shady past and is not as perfect as he appears. Thriller, starring Josie Davis and Marc Menard.(n)
Channel 5|1464105600|5 News at 5|24/05/2016||0|0|News|Sian Williams presents a round-up of the day's headlines from around the world.(n)
Channel 5|1464107400|Neighbours|||0|0|Soap,Melodrama|Brodie divulges a piece of detail regarding the Lassiter's blast that he should not know. Terese seeks distraction from her grief, while Lauren feels uneasy about Ned.(n)
Channel 5|1464109200|Home and Away|||0|0|Soap,Melodrama|Zac is forced to perform life-saving emergency surgery on Hunter, Skye teases VJ when she realises he has a crush on Billie, and Greg finds out Zac was in prison with his son Wayne.(n)
Channel 5|1464111000|5 News Tonight|24/05/2016||0|0|General News,Current Affairs|A round-up of the evening's headlines, including coverage of the latest national and international stories.(n)
Channel 5|1464112500|Referendum Campaign Broadcast|||0|0|General Social,Political Issues,Economics|By the Britain Stronger in Europe campaign.(n)
Channel 5|1464112800|FIA World Rally Championship Highlights|2016 Rally de Portugal||1|5|Rallying|The Rally de Portugal. Jon Desborough presents highlights of the fifth round of the season, based in the northern city and municipality of Matosinhos. This round was set to feature a total of 19 stages covering 368km, all of which featured gravel roads.(n)
Channel 5|1464116400|The Yorkshire Vet|||2|7|General Arts,Culture|Julian Norton and his practice partner Peter Wright have to cope with night-time emergencies, as Julian performs outdoor surgery on a first-time mum and Peter examines a cat with a potentially life-threatening condition. Newly qualified vet Esme Telfer performs her first emergency caesarian at the Skeldale practice, while at Green's farm Treacle the calf falls ill and it is touch-and-go whether she will survive. Later, a pack of bloodhound pups causes chaos in the surgery.(n)
Channel 5|1464120000|The KKK: Behind The Mask|||0|0|General Education,Science|The Ku Klux Klan is the most notorious white supremacist group in America. Once having over a million members, today it's a shadow of its former self, and yet the marches, the cross burnings and the racial hatred continues in the Southern states. This documentary profiles today's Klan members, examines the impact the group has had on America over the last 150 years, and examines whether America is heading for a new race war.(n)
Channel 5|1464123600|Your Child In Their Hands|Your Child In Their Hands: Kids' Hospital||1|2|General Arts,Culture|The documentary exploring the trials faced by families at Royal Manchester Children's Hospital continues, as parents-to-be Lizzie and her partner Andy come to terms with the fact that their unborn baby will need urgent treatment to survive. Teenager Connor discovers he has a very rare condition that causes his immune system to attack his own body, and the news proves devastating for his father Ian, whose family has been hit by tragedy two times before. Plus, a youngster drifting in and out of consciousness provides cause for concert for A&E staff, and a mother's concerns get the better of her as her son goes into theatre for an operation on his leg.(n)
Channel 5|1464127200|Up Late with Rylan|||1|10|Talk Show|Rylan Clark-Neal hosts the chat show, featuring celebrity guests and music as well as games for the studio audience and the viewers at home.(n)
Channel 5|1464129900|Can't Pay? We'll Take It Away|||4|6|Documentary|Agents Stewart and Vic experience one of the most violent cases they have ever faced when they are confronted by an angry older gentleman. Later, the pair chase £3,000 owed for an unwanted car engine, but the debtor is convinced that he knows the law and the agents' jobs better than they do. Meanwhile, Steve and Ben face a dilemma in north London, where a tenant is being evicted for rent arrears, and in south London, Paul and Steve have no option but to force a dramatic entry into a property.(n)
Sky Sports 1|1463877000|Barclays Premier League Legends|PL Legends: Alan Shearer||0|0|Football - Club|A profile of former Newcastle United, Blackburn Rovers and England striker Alan Shearer.
Sky Sports 1|1463878800|Football Gold|Manchester United v Liverpool: 2013/14||0|0|Football,Soccer|Manchester United v Liverpool from the 2013/14 Premier League season.
Sky Sports 1|1463879700|Football Gold|Tottenham Hotspur v Arsenal: 2013/14||0|0|Football,Soccer|Tottenham Hotspur v Arsenal from the 2013/14 Premier League season.
Sky Sports 1|1463880600|Football Gold|Sunderland v West Ham United: 2013/14||0|0|Football,Soccer|Sunderland v West Ham United from the 2013/14 Premier League season.
Sky Sports 1|1463881500|Football Gold|Tottenham Hotspur v Liverpool: 2013/14||0|0|Football,Soccer|Tottenham Hotspur v Liverpool from the 2013/14 Premier League season.
Sky Sports 1|1463882400|Barclays Premier League Legends|PL Legends: Robbie Fowler||0|0|Football - Club|A look back at the career of striker Robbie Fowler who scored 162 Premier League goals during spells with Liverpool, Manchester City, Leeds United and Blackburn Rovers.
Sky Sports 1|1463884200|Premier League Years|1992/93||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 1992/93 season, all set to a specially selected soundtrack from the time.
Sky Sports 1|1463891400|Football Gold|Manchester United v Liverpool: 2013/14||0|0|Football,Soccer|Manchester United v Liverpool from the 2013/14 Premier League season.
Sky Sports 1|1463892300|Football Gold|Tottenham Hotspur v Arsenal: 2013/14||0|0|Football,Soccer|Tottenham Hotspur v Arsenal from the 2013/14 Premier League season.
Sky Sports 1|1463893200|Football Gold|Chelsea v Tottenham Hotspur: 1993/94||0|0|Football,Soccer|Classic archive action from 1993/94 when Chelsea met Tottenham Hotspur at Stamford Bridge.
Sky Sports 1|1463894100|Football Gold|Arsenal v Leeds United: 2002/03||0|0|Football,Soccer|Action from the Premiership clash between Arsenal and Leeds United in the 2002/03 season.
Sky Sports 1|1463895000|Football Gold|West Ham United v Tottenham Hotspur: 2006/07||0|0|Football,Soccer|West Ham United v Tottenham Hotspur. A chance to relive the classic Premier League encounter from the 2006/07 season.
Sky Sports 1|1463895900|Football Gold|Manchester City v Tottenham Hotspur: 2002/03||0|0|Football,Soccer|Manchester City v Tottenham Hotspur. Classic archive action from the 2002/03 clash between the sides.
Sky Sports 1|1463896800|Barclays Premier League Legends|PL Legends: Juninho||0|0|Football - Club|A profile of Middlesbrough's former Brazilian midfielder Juninho.
Sky Sports 1|1463898600|Premier League 100 Club|PL 100 Club: Ian Wright||0|0|Football - Club|A look at Ian Wright's top-flight goals.
Sky Sports 1|1463900400|Scottish Cup Football|Rangers v Hibernian||0|0|Football - Club|Rangers v Hibernian. Action from the final at Hampden Park, which was the first-ever to be contested between two clubs from the second tier.
Sky Sports 1|1463904000|Live HSBC Sevens World Series|2015/16 London Sevens: Day Two Session One||0|0|Rugby Union - International|The London Sevens. Coverage of day two of the 10th and final round of the season, which comes from Twickenham.
Sky Sports 1|1463916600|Live First Utility Super League|Live Super League Magic Weekend: Wakefield Trinity Wildcats v Catalan Dragons||0|0|Rugby League - Domestic|Wakefield Trinity Wildcats v Catalan Dragons (Kick-off 1.00pm). Coverage of the match from St James' Park in Newcastle, as the 15th round of fixtures continues on Magic Weekend.
Sky Sports 1|1463925600|Live First Utility Super League|Live Super League Magic Weekend: St Helens v Huddersfield Giants||0|0|Rugby League - Domestic|St Helens v Huddersfield Giants (Kick-off 3.15pm). Coverage of the match from St James' Park in Newcastle, as the 15th round of fixtures continues on Magic Weekend.
Sky Sports 1|1463933700|Live First Utility Super League|Live Super League Magic Weekend: Hull FC v Hull Kingston Rovers||0|0|Rugby League - Domestic|Hull FC v Hull Kingston Rovers (Kick-off 5.30pm). Coverage of the match from St James' Park in Newcastle, as the 15th round of fixtures concludes on Magic Weekend. The most recent meeting between the sides saw FC come back from 20-0 down with just quarter of the match remaining to record a remarkable 22-20 victory at Craven Park on Good Friday.
Sky Sports 1|1463943600|Live Copa Del Rey Football|Live Copa Del Rey Final: Barcelona v Sevilla||0|0|Football,Soccer|Barcelona v Sevilla (Kick-off 8.30pm). Coverage of the showpiece match from Estadio Vicente Calderon in Madrid.(c)
Sky Sports 1|1463954400|Scottish Cup Football|Rangers v Hibernian||0|0|Football - Club|Rangers v Hibernian. Action from the final at Hampden Park, which was the first-ever to be contested between two clubs from the second tier.(c)
Sky Sports 1|1463958000|Copa Del Rey Football|Barcelona v Sevilla||0|0|Football - Club|Barcelona v Sevilla. Action from the final of the showpiece occasion in Spanish cup football, which took place at the Vicente Calderon.(c)
Sky Sports 1|1463958900|Live MLS|Los Angeles Galaxy v San Jose Earthquakes||0|0|Football - Club|Los Angeles Galaxy v San Jose Earthquakes (Kick-off TBA). Coverage of the Western Conference clash from StubHub Centre.(c)
Sky Sports 1|1463966700|My Greatest Game|Martin Tyler||0|0|Football,Soccer|Martin Tyler discusses Liverpool v Newcastle United from April 1996.(c)
Sky Sports 1|1463967000|Football Gold|Chelsea v Manchester City 2009/10||0|0|Football,Soccer|Action from the Premier League match between Chelsea and Manchester City in the 2009/10 season.
Sky Sports 1|1463967900|Football Gold|Manchester City v Manchester United: 1993/94||0|0|Football,Soccer|A look back at the Premiership match between Manchester City and Manchester United from the 1993/94 season.
Sky Sports 1|1463968800|Barclays Premier League Legends|PL Legends: Paolo Di Canio||0|0|Football - Club|A profile of Paolo Di Canio, the former Sheffield Wednesday, West Ham United and Charlton Athletic forward who scored 67 goals in almost 200 Premier League appearances.
Sky Sports 1|1463970600|Premier League 100 Club|PL 100 Club: Frank Lampard||0|0|Football - Club|A chance to relive the goals of Frank Lampard, who scored more than any other midfielder in Premier League history during his time with West Ham United, Chelsea and Manchester City.
Sky Sports 1|1463972400|Premier League Years|1994/95||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 1994/95 season, all set to a specially selected soundtrack from the time.
Sky Sports 1|1463979600|Football Gold|Chelsea v Manchester United: 2013/14||0|0|Football,Soccer|Chelsea v Manchester United. Highlights of the Premier League clash from the 2013/14 season, which came from Stamford Bridge.
Sky Sports 1|1463980500|Football Gold|Aston Villa v West Bromwich Albion: 2013/14||0|0|Football,Soccer|Aston Villa v West Bromwich Albion. Action from the 2013/14 Premier League clash at Villa Park.
Sky Sports 1|1463981400|Football Gold|Chelsea v Manchester City 2009/10||0|0|Football,Soccer|Action from the Premier League match between Chelsea and Manchester City in the 2009/10 season.
Sky Sports 1|1463982300|Football Gold|Manchester United v Arsenal: 2011/12||0|0|Football,Soccer|A chance to relive the Premier League contest between Manchester United and Arsenal at Old Trafford from August 2011.
Sky Sports 1|1463983200|WWE: Raw|||0|0|Wrestling|Wrestling action from the States with the over-the-top stars, featuring the likes of Randy Orton and John Cena. Presented by Michael Cole, John `Bradshaw' Layfield and Byron Saxton.
Sky Sports 1|1463986800|Premier League 100 Club|PL 100 Club: Didier Drogba||0|0|Football - Club|The best of Didier Drogba's 104 Premier League goals for Chelsea, which were scored over two spells with the club between 2004 and 2015.
Sky Sports 1|1463988600|Barclays Premier League Legends|PL Legends: Gianfranco Zola||0|0|Football - Club|A profile of former Chelsea forward Gianfranco Zola.
Sky Sports 1|1463990400|Major League Soccer|MLS Highlights: Portland Timbers v Vancouver Whitecaps||0|0|Football - Club|Portland Timbers v Vancouver Whitecaps. Action from the Western Conference clash at Providence Park.
Sky Sports 1|1463997600|Major League Soccer|MLS Highlights: Los Angeles Galaxy v San Jose Earthquakes||0|0|Football - Club|Los Angeles Galaxy v San Jose Earthquakes. Action from the Western Conference clash at StubHub Centre.
Sky Sports 1|1464004800|Premier League Years|1993/94||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 1993/94 season, all set to a specially selected soundtrack from the time.
Sky Sports 1|1464012000|Scottish Cup Football|Rangers v Hibernian||0|0|Football - Club|Rangers v Hibernian. Action from the final at Hampden Park, which was the first-ever to be contested between two clubs from the second tier.
Sky Sports 1|1464015600|Copa Del Rey Football|Barcelona v Sevilla||0|0|Football - Club|Barcelona v Sevilla. Action from the final of the showpiece occasion in Spanish cup football, which took place at the Vicente Calderon.
Sky Sports 1|1464016500|Football Gold|Aston Villa v West Bromwich Albion: 2013/14||0|0|Football,Soccer|Aston Villa v West Bromwich Albion. Action from the 2013/14 Premier League clash at Villa Park.
Sky Sports 1|1464017400|Football Gold|Chelsea v Manchester City 2009/10||0|0|Football,Soccer|Action from the Premier League match between Chelsea and Manchester City in the 2009/10 season.
Sky Sports 1|1464018300|Football Gold|Manchester United v Arsenal: 2011/12||0|0|Football,Soccer|A chance to relive the Premier League contest between Manchester United and Arsenal at Old Trafford from August 2011.
Sky Sports 1|1464019200|Football's Greatest Players|Michael Laudrup||0|0|Football - International|The career of former Barcelona, Real Madrid and Denmark star Michael Laudrup. The attacking midfielder won many honours during his career, including four La Liga titles with Barcelona and one with Real Madrid, and also represented his country on 104 occasions.
Sky Sports 1|1464021000|Fantasy Football Club - The Highlights|2015/16||0|0|Football - Club|Max Rushden and Paul Merson look back on highlights of the show, which focusses on key fantasy football issues, and features studio guests.
Sky Sports 1|1464022800|Scottish Cup Football|Rangers v Hibernian||0|0|Football - Club|Rangers v Hibernian. Action from the final at Hampden Park, which was the first-ever to be contested between two clubs from the second tier.
Sky Sports 1|1464026400|Football Gold|Aston Villa v West Bromwich Albion: 2013/14||0|0|Football,Soccer|Aston Villa v West Bromwich Albion. Action from the 2013/14 Premier League clash at Villa Park.
Sky Sports 1|1464027300|Copa Del Rey Football|Barcelona v Sevilla||0|0|Football - Club|Barcelona v Sevilla. Action from the final of the showpiece occasion in Spanish cup football, which took place at the Vicente Calderon.
Sky Sports 1|1464028200|Live Elite League Speedway|Poole Pirates v Belle Vue Aces||0|0|Motorcycling|Poole Pirates v Belle Vue Aces. Coverage of the top-flight meeting at Poole Stadium.
Sky Sports 1|1464035400|First Utility Super League Highlights|Magic Weekend Highlights: Salford Red Devils v Widnes Vikings||0|0|Rugby League - Domestic|Salford Red Devils v Widnes Vikings. Action from the Super League match at St James' Park in Newcastle.
Sky Sports 1|1464036300|First Utility Super League Highlights|Magic Weekend Highlights: Warrington Wolves v Castleford Tigers||0|0|Rugby League - Domestic|Warrington Wolves v Castleford Tigers. Action from the Super League match at St James' Park in Newcastle.
Sky Sports 1|1464037200|First Utility Super League Highlights|Magic Weekend Highlights: Leeds Rhinos v Wigan Warriors||0|0|Rugby League - Domestic|Leeds Rhinos v Wigan Warriors. Action from the Super League match at St James' Park in Newcastle.
Sky Sports 1|1464038100|First Utility Super League Highlights|Magic Weekend Highlights: Wakefield Trinity Wildcats v Catalan Dragons||0|0|Rugby League - Domestic|Wakefield Trinity Wildcats v Catalan Dragons. Action from the Super League match at St James' Park in Newcastle.
Sky Sports 1|1464039000|First Utility Super League Highlights|Magic Weekend Highlights: St Helens v Huddersfield Giants||0|0|Rugby League - Domestic|St Helens v Huddersfield Giants. Action from the Super League match at St James' Park in Newcastle.
Sky Sports 1|1464039900|First Utility Super League Highlights|Magic Weekend Highlights: Hull FC v Hull Kingston Rovers||0|0|Rugby League - Domestic|Hull FC v Hull Kingston Rovers. Action from the Super League match at St James' Park in Newcastle.
Sky Sports 1|1464040800|Elite League Speedway|Poole Pirates v Belle Vue Aces||0|0|Motorcycling|Poole Pirates v Belle Vue Aces. Action from the top-flight meeting at Poole Stadium.
Sky Sports 1|1464048000|First Utility Super League Highlights|Magic Weekend Highlights: Salford Red Devils v Widnes Vikings||0|0|Rugby League - Domestic|Salford Red Devils v Widnes Vikings. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 1|1464048900|First Utility Super League Highlights|Magic Weekend Highlights: Warrington Wolves v Castleford Tigers||0|0|Rugby League - Domestic|Warrington Wolves v Castleford Tigers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 1|1464049800|First Utility Super League Highlights|Magic Weekend Highlights: Leeds Rhinos v Wigan Warriors||0|0|Rugby League - Domestic|Leeds Rhinos v Wigan Warriors. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 1|1464050700|First Utility Super League Highlights|Magic Weekend Highlights: Wakefield Trinity Wildcats v Catalan Dragons||0|0|Rugby League - Domestic|Wakefield Trinity Wildcats v Catalan Dragons. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 1|1464051600|First Utility Super League Highlights|Magic Weekend Highlights: St Helens v Huddersfield Giants||0|0|Rugby League - Domestic|St Helens v Huddersfield Giants. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 1|1464052500|First Utility Super League Highlights|Magic Weekend Highlights: Hull FC v Hull Kingston Rovers||0|0|Rugby League - Domestic|Hull FC v Hull Kingston Rovers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 1|1464053400|Premier League Years|2008/09||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 2008/09 season, all set to a specially selected soundtrack from the time.(n)
Sky Sports 1|1464060600|Barclays Premier League Legends|PL Legends: David Seaman||0|0|Football - Club|The career of David Seaman, who was Arsenal's number one goalkeeper for the first 11 seasons of the Premier League, before moving to Manchester City in 2003 and retiring in 2004.(n)
Sky Sports 1|1464062400|Premier League 100 Club|PL 100 Club: Emile Heskey||0|0|Football - Club|The best of Emile Heskey's top-flight goals, which he scored with five different clubs - Leicester City, Liverpool, Birmingham City, Wigan Athletic and Aston Villa.(n)
Sky Sports 1|1464064200|Premier League 100 Club|PL 100 Club: Frank Lampard||0|0|Football - Club|A chance to relive the goals of Frank Lampard, who scored more than any other midfielder in Premier League history during his time with West Ham United, Chelsea and Manchester City.(n)
Sky Sports 1|1464066000|Football Gold|Everton v Manchester City: 2013/14||0|0|Football,Soccer|Everton v Manchester City. Action from the top-flight match at Goodison Park from the 2013/14 season.(n)
Sky Sports 1|1464066900|Football Gold|Chelsea v Manchester United: 2011/12||0|0|Football,Soccer|Chelsea v Manchester United. Highlights of the Premier League clash from the 2011/12 season, which came from Stamford Bridge and ended in a 3-3 draw.(n)
Sky Sports 1|1464067800|Football Gold|Cardiff City v Liverpool: 2013/14||0|0|Football,Soccer|Cardiff City v Liverpool from the 2013/14 Premier League season.(n)
Sky Sports 1|1464068700|Football Gold|West Bromwich Albion v Cardiff City: 2013/14||0|0|Football,Soccer|West Bromwich Albion v Cardiff City. A chance to relive the classic 2013/14 Premier League match from the Hawthorns.(n)
Sky Sports 1|1464069600|WWE: Smackdown|||0|0|Wrestling|Spectacular grappling action with the over-the-top stars of the States, profiling fighters causing a stir and following feuds as they spill out of the ring.(n)
Sky Sports 1|1464073200|Premier League 100 Club|PL 100 Club: Steven Gerrard||0|0|Football - Club|A chance to relive the league goals scored by Steven Gerrard. The influential former Liverpool captain is the second-highest-scoring midfielder in Premier League history with 120.(n)
Sky Sports 1|1464075000|Barclays Premier League Legends|PL Legends: Jamie Carragher||0|0|Football - Club|The career of former Liverpool defender Jamie Carragher, who made 508 Premier League appearances for his home town club between 1997 and 2013.(n)
Sky Sports 1|1464076800|Premier League Years|2001/02||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 2001/02 season, all set to a specially selected soundtrack from the time.(n)
Sky Sports 1|1464084000|Fantasy Football Club - The Highlights|2015/16||0|0|Football - Club|Max Rushden and Paul Merson look back on highlights of the show, which focusses on key fantasy football issues, and features studio guests.(n)
Sky Sports 1|1464085800|Football Gold|Cardiff City v Liverpool: 2013/14||0|0|Football,Soccer|Cardiff City v Liverpool from the 2013/14 Premier League season.(n)
Sky Sports 1|1464086700|Football Gold|West Bromwich Albion v Cardiff City: 2013/14||0|0|Football,Soccer|West Bromwich Albion v Cardiff City. A chance to relive the classic 2013/14 Premier League match from the Hawthorns.(n)
Sky Sports 1|1464087600|Premier League 100 Club|PL 100 Club: Frank Lampard||0|0|Football - Club|A chance to relive the goals of Frank Lampard, who scored more than any other midfielder in Premier League history during his time with West Ham United, Chelsea and Manchester City.(n)
Sky Sports 1|1464089400|Barclays Premier League Legends|PL Legends: Paolo Di Canio||0|0|Football - Club|A profile of Paolo Di Canio, the former Sheffield Wednesday, West Ham United and Charlton Athletic forward who scored 67 goals in almost 200 Premier League appearances.(n)
Sky Sports 1|1464091200|Premier League Years|1994/95||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 1994/95 season, all set to a specially selected soundtrack from the time.(n)
Sky Sports 1|1464098400|Live Indian Premier League|2016 Qualifying Play-Off One||0|0|Cricket - Domestic|Coverage of the first qualifying play-off match from M Chinnaswamy Stadium in Bangalore, where two teams compete for a place in the final.(n)
Sky Sports 1|1464114600|Cricket Classics|England v Australia: Second Test 2005||0|0|Cricket - Domestic|England v Australia. Highlights of the Second Ashes Test at Edgbaston from 2005.(n)
Sky Sports 1|1464115500|Cricket Classics|South Africa v Australia: Fifth ODI 2006||0|0|Cricket - Domestic|South Africa v Australia. Action from the fifth one-day international between the sides at New Wanderers Stadium, Johannesburg in 2006.(n)
Sky Sports 1|1464116400|Indian Premier League|2016 Qualifying Play-Off One||0|0|Cricket - Domestic|Action from the first qualifying play-off match at M Chinnaswamy Stadium in Bangalore, where two teams competed for a place in the final.(n)
Sky Sports 2|1463871600|Cricket's Greatest|Wasim Akram||0|0|Cricket - International|A profile of former Pakistan fast bowler Wasim Akram.
Sky Sports 2|1463873400|Live MLS|Orlando City SC v Montreal Impact||0|0|Football - Club|Orlando City SC v Montreal Impact (Kick-off 12.30am). Coverage of the Eastern Conference match from Orlando Citrus Bowl in Florida.
Sky Sports 2|1463880600|Test Cricket|England v Sri Lanka: First Test Day Three||0|0|Cricket - International|England v Sri Lanka. Highlights of the third day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1463884200|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Three||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the third day of the First Test at Headingley.
Sky Sports 2|1463887800|Cricket's Greatest|Graeme Pollock||0|0|Cricket - International|A profile of former South Africa batsman Graeme Pollock.
Sky Sports 2|1463889600|Cricket Classics|West Indies v South Africa: 2005 ODI||0|0|Cricket - Domestic|Action from the third one-dayer between West Indies and South Africa from 2005, held at Kingston Oval in Bridgetown, Barbados.
Sky Sports 2|1463893200|Indian Premier League|Rising Pune Supergiants v Kings XI Punjab||0|0|Cricket - Domestic|Rising Pune Supergiants v Kings XI Punjab. Highlights of the match from the Twenty20 competition, held at Maharashtra Cricket Association Stadium in Pune.
Sky Sports 2|1463896800|Indian Premier League|Gujarat Lions v Mumbai Indians||0|0|Cricket - Domestic|Gujarat Lions v Mumbai Indians. Action from the Twenty20 match, which took place at Green Park in Kanpur.
Sky Sports 2|1463900400|Test Cricket|England v Sri Lanka: First Test Day Three||0|0|Cricket - International|England v Sri Lanka. Highlights of the third day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1463904000|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Three||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the third day of the First Test at Headingley.
Sky Sports 2|1463907600|Cricket Writers on TV|22 May 2016||0|0|Cricket - International|Paul Allott is joined by a trio of cricket journalists to discuss the latest issues making waves in the sport over the past seven days.
Sky Sports 2|1463909400|Live Test Cricket|England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. Coverage of the fourth day of the First Test at Headingley, where the three-match series continues.
Sky Sports 2|1463940000|Cricket in the 90s|Cricket in the 90s - England in the 90s||0|0|Cricket - International|Documentary looking back at the national team's performances in the decade.
Sky Sports 2|1463943600|Test Cricket|England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. Highlights of the fourth day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1463947200|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fourth day of the First Test at Headingley.
Sky Sports 2|1463950800|Indian Premier League|Kolkata Knight Riders v Sunrisers Hyderabad||0|0|Cricket - Domestic|Kolkata Knight Riders v Sunrisers Hyderabad. A chance to see the Twenty20 encounter at Eden Gardens, where the lucrative competition continued.
Sky Sports 2|1463954400|Indian Premier League|Delhi Daredevils v Royal Challengers Bangalore||0|0|Cricket - Domestic|Delhi Daredevils v Royal Challengers Bangalore. Action from the group-stage match in the Twenty20 competition, from Feroz Shah Kotla.
Sky Sports 2|1463958000|Cricket Classics|England v Australia: 2005 Natwest Series Game Three||0|0|Cricket - Domestic|England v Australia. Action from match three of the 2005 Natwest Series, held at the County Ground in Bristol.
Sky Sports 2|1463958900|Cricket Classics|England v Australia: 2005 Natwest Final||0|0|Cricket - Domestic|Highlights of the 2005 Natwest series final between England and Australia, which was held at Lord's.
Sky Sports 2|1463959800|Cricket's Greatest|Sachin Tendulkar||0|0|Cricket - International|A profile of Sachin Tendulkar, regarded as one of the most outstanding talents ever to play the sport.
Sky Sports 2|1463961600|Test Cricket|England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. Highlights of the fourth day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1463965200|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fourth day of the First Test at Headingley.
Sky Sports 2|1463968800|Cricket Classics|England v India: 2002 Natwest Series Final||0|0|Cricket - Domestic|England v India in the 2002 Natwest Series final.
Sky Sports 2|1463969700|Cricket Classics|England v Australia: Second Test 2005||0|0|Cricket - Domestic|England v Australia. Highlights of the Second Ashes Test at Edgbaston from 2005.
Sky Sports 2|1463970600|Cricket's Greatest|Sunil Gavaskar||0|0|Cricket - International|A profile of Sunil Gavaskar, the former Indian opening batsman, whose run-scoring was prolific at the top of the order.
Sky Sports 2|1463972400|Test Cricket|England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. Highlights of the fourth day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1463976000|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fourth day of the First Test at Headingley.
Sky Sports 2|1463979600|Cricket's Greatest|Don Bradman||0|0|Cricket - International|A profile of Don Bradman.
Sky Sports 2|1463981400|Cricket's Greatest|Garfield Sobers||0|0|Cricket - International|A profile of Garfield Sobers.
Sky Sports 2|1463983200|Test Cricket|England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. Highlights of the fourth day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1463986800|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Four||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fourth day of the First Test at Headingley.
Sky Sports 2|1463990400|Cricket's Greatest|Wasim Akram||0|0|Cricket - International|A profile of former Pakistan fast bowler Wasim Akram.
Sky Sports 2|1463992200|Cricket's Greatest|Graeme Pollock||0|0|Cricket - International|A profile of former South Africa batsman Graeme Pollock.
Sky Sports 2|1463994000|AB de Villiers Masterclass|||0|0|Cricket - International|A cricketing masterclass with the South Africa captain.
Sky Sports 2|1463995800|Live Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Coverage of the fifth and final day of the First Test at Headingley, where the three-match series continues.
Sky Sports 2|1464022800|Cricket's Greatest|Ian Botham||0|0|Cricket - International|A profile of former England cricketer Ian Botham, regarded as one of the greatest all-rounders in the history of the sport.
Sky Sports 2|1464024600|Cricket's Greatest|Graham Gooch||0|0|Cricket - International|A profile of former England batsman Graham Gooch, who remains one of the leading run-scorers for his country following a long and successful career as an opener.
Sky Sports 2|1464026400|Sporting Heroes|Sporting Heroes: Peter Schmeichel Interviews Peter Shilton||0|0|General Sports|A conversation between the two former goalkeepers, who are ranked among the best of all time.
Sky Sports 2|1464030000|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1464033600|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.
Sky Sports 2|1464037200|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.
Sky Sports 2|1464040800|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.
Sky Sports 2|1464044400|Cricket Classics|England v Australia: 2005 Natwest Final||0|0|Cricket - Domestic|Highlights of the 2005 Natwest series final between England and Australia, which was held at Lord's.(n)
Sky Sports 2|1464048000|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.(n)
Sky Sports 2|1464051600|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.(n)
Sky Sports 2|1464055200|Cricket's Greatest|Steve Waugh||0|0|Cricket - International|A profile of former Australia captain Steve Waugh, regarded as one of the greatest all-rounders and leaders in the sport's modern history.(n)
Sky Sports 2|1464057000|Cricket's Greatest|Dennis Lillee||0|0|Cricket - International|A profile of Dennis Lillee, one of the most feared fast bowlers in the history of the sport.(n)
Sky Sports 2|1464058800|Cricket's Greatest|Allan Border||0|0|Cricket - International|A profile of Allan Border, the former Australian captain, who helped to turn his nation's fortunes around in the late 1980s.(n)
Sky Sports 2|1464060600|Cricket's Greatest|Glenn McGrath||0|0|Cricket - International|A profile of former Australia bowler Glenn McGrath.(n)
Sky Sports 2|1464062400|Time of Our Lives|Olympics Munich 1972||0|0|General Sports|Mary Peters, Mark Phillips and Rodney Pattisson look back at their gold medal-winning performances for Great Britain at the 1972 Munich Olympics, in athletics' pentathlon, equestrian's three-day event team competition and sailing respectively.(n)
Sky Sports 2|1464066000|Cricket's Greatest|Ian Botham||0|0|Cricket - International|A profile of former England cricketer Ian Botham, regarded as one of the greatest all-rounders in the history of the sport.(n)
Sky Sports 2|1464067800|Cricket's Greatest|David Gower||0|0|Cricket - International|A profile of former England batsman David Gower, who was one of the leading players in the sport during the 1980s, and became known for his flamboyant stroke making.(n)
Sky Sports 2|1464069600|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.(n)
Sky Sports 2|1464073200|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.(n)
Sky Sports 2|1464076800|First Utility Super League Highlights|Magic Weekend Highlights: Salford Red Devils v Widnes Vikings||0|0|Rugby League - Domestic|Salford Red Devils v Widnes Vikings. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 2|1464077700|First Utility Super League Highlights|Magic Weekend Highlights: Warrington Wolves v Castleford Tigers||0|0|Rugby League - Domestic|Warrington Wolves v Castleford Tigers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 2|1464078600|First Utility Super League Highlights|Magic Weekend Highlights: Leeds Rhinos v Wigan Warriors||0|0|Rugby League - Domestic|Leeds Rhinos v Wigan Warriors. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 2|1464079500|First Utility Super League Highlights|Magic Weekend Highlights: Wakefield Trinity Wildcats v Catalan Dragons||0|0|Rugby League - Domestic|Wakefield Trinity Wildcats v Catalan Dragons. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 2|1464080400|First Utility Super League Highlights|Magic Weekend Highlights: St Helens v Huddersfield Giants||0|0|Rugby League - Domestic|St Helens v Huddersfield Giants. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 2|1464081300|First Utility Super League Highlights|Magic Weekend Highlights: Hull FC v Hull Kingston Rovers||0|0|Rugby League - Domestic|Hull FC v Hull Kingston Rovers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 2|1464082200|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.(n)
Sky Sports 2|1464085800|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.(n)
Sky Sports 2|1464089400|Cricket's Greatest|Ian Botham||0|0|Cricket - International|A profile of former England cricketer Ian Botham, regarded as one of the greatest all-rounders in the history of the sport.(n)
Sky Sports 2|1464091200|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.(n)
Sky Sports 2|1464094800|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.(n)
Sky Sports 2|1464098400|Barclays Premier League Legends|PL Legends: Juninho||0|0|Football - Club|A profile of Middlesbrough's former Brazilian midfielder Juninho.(n)
Sky Sports 2|1464100200|Premier League 100 Club|PL 100 Club: Teddy Sheringham||0|0|Football - Club|The best of Teddy Sheringham's 146 Premier League goals scored with five different clubs - Nottingham Forest, Tottenham Hotspur, Manchester United, Portsmouth and West Ham United.(n)
Sky Sports 2|1464102000|Test Cricket|England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. Highlights of the fifth and final day of the First Test at Headingley, where the three-match series continued.(n)
Sky Sports 2|1464105600|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Five||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the fifth and final day of the First Test at Headingley.(n)
Sky Sports 2|1464109200|Premier League 100 Club|PL 100 Club: Andy Cole||0|0|Football - Club|The best of Andy Cole's 187 goals in the Premier League, scored for Newcastle United, Manchester United, Blackburn Rovers, Manchester City, Fulham, Portsmouth and Birmingham City.(n)
Sky Sports 2|1464111000|Premier League 100 Club|PL 100 Club: Dwight Yorke||0|0|Football - Club|A chance to relive the best of Dwight Yorke's 123 goals in the Premier League, which he scored for Aston Villa, Manchester United, Blackburn Rovers, Birmingham City and Sunderland.(n)
Sky Sports 2|1464112800|Live Greyhound Racing|2016 William Hill Derby Quarter-Finals||0|0|Greyhound Racing|Coverage of this evening's William Hill Derby quarter-finals at Wimbledon, where the top three in each race will book their place in the semi-finals.(n)
Sky Sports 2|1464121800|Sky Sports Boxing Gold|Carl Froch v Lucian Bute||0|0|Boxing|Lucian Bute v Carl Froch. Action from the 2012 bout for the IBF Super Middleweight title at the Nottingham Arena, where Bute was making the 10th defence of his title.(n)
Sky Sports 2|1464123600|Cricket's Greatest|Shane Warne||0|0|Cricket - International|A profile of Shane Warne, who is widely regarded as one of the greatest spin bowlers of all time.(n)
Sky Sports 2|1464125400|MLS Round-Up Show|2016||0|0|Football - Club|A review of the latest round of Major League Soccer fixtures.(n)
Sky Sports 2|1464127200|Time of Our Lives|The Ramsey Years||0|0|General Sports|Ray Crawford, Ted Phillips and Larry Carberry join Jeff Stelling to reminisce about Ipswich Town's incredible season of 1961/62, which saw them win the league and face the likes of Fiorentina and AC Milan in the European Cup.(n)
Sky Sports 3|1463873400|The Verdict|Test Cricket: The Verdict: England v Sri Lanka: First Test Day Three||0|0|Cricket - International|England v Sri Lanka. A panel of guests discuss the third day of the First Test at Headingley.
Sky Sports 3|1463877000|Sporting Triumphs|Jamie Carragher Winning 2005 Champions League||0|0|General Sports|Jamie Carragher relives Liverpool's dramatic 2005 Champions League final victory over AC Milan, when they came back from 3-0 down to eventually win 3-2 on penalties.
Sky Sports 3|1463877900|Sporting Triumphs|Sean Fitzpatrick - All Blacks Win First Rugby World Cup||0|0|General Sports|Former All Black Sean Fitzpatrick takes a look back at how New Zealand won the inaugural Rugby World Cup in 1987, which was staged in Australia and New Zealand.
Sky Sports 3|1463878800|Sky Sports Boxing Gold|Carl Froch v Lucian Bute||0|0|Boxing|Lucian Bute v Carl Froch. Action from the 2012 bout for the IBF Super Middleweight title at the Nottingham Arena, where Bute was making the 10th defence of his title.
Sky Sports 3|1463880600|Fight Night International|Joseph Parker v Carlos Takam||0|0|Boxing|Joseph Parker v Carlos Takam. Action from the heavyweight bout, a final eliminator for Anthony Joshua's IBF world title that took place at the Vodafone Events Centre in Auckland.
Sky Sports 3|1463887800|Sporting Greats|Seve Ballesteros||0|0|General Sports|A profile of Seve Ballesteros, who won five golf Majors and tasted Ryder Cup glory four times as a player and on another occasion as a team captain. The Spaniard gained many admirers due to his flamboyant style of play before dying of brain cancer in May 2011.
Sky Sports 3|1463889600|Darts Gold|WDC Finals 06/07||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2006 and 2007.
Sky Sports 3|1463891400|Darts Gold|WDC Finals 08/09||0|0|Darts|Action from the 2008 and 2009 World Darts Championship finals.
Sky Sports 3|1463893200|Darts Gold|WDC Finals 10/11||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2010 and 2011.
Sky Sports 3|1463895000|Darts Gold|WDC Finals 12/13||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2012 and 2013.
Sky Sports 3|1463896800|Time of Our Lives|Champion Jockeys||0|0|General Sports|Former jockeys Willie Carson, Pat Eddery and Joe Mercer look back on their careers.
Sky Sports 3|1463900400|Major League Soccer|MLS Highlights: Chicago Fire v Houston Dynamo||0|0|Football - Club|Chicago Fire v Houston Dynamo. Action from the top-flight encounter at Toyota Park.
Sky Sports 3|1463907600|Major League Soccer|MLS Highlights: New York City FC v New York Red Bulls||0|0|Football - Club|New York City FC v New York Red Bulls. Action from the Eastern Conference match, which was held at Yankee Stadium.
Sky Sports 3|1463914800|Barclays Premier League Legends|PL Legends: Alan Shearer||0|0|Football - Club|A profile of former Newcastle United, Blackburn Rovers and England striker Alan Shearer.
Sky Sports 3|1463916600|Live HSBC Sevens World Series|2016 London Sevens: Day Two||0|0|Rugby Union - International|The London Sevens. Coverage of the second and concluding day of the 10th and final round of the season, which takes place at Twickenham. The climax of the season at the home of English rugby will see the successor being crowned to last year's winners FIji.
Sky Sports 3|1463940000|Super Rugby Try Time|2016||0|0|Rugby League - Domestic|A round-up of all the tries, highlights and news headlines from the most recent round of the Super Rugby season.
Sky Sports 3|1463941800|Major League Soccer|MLS Highlights: Orlando City SC v Montreal Impact||0|0|Football - Club|Orlando City SC v Montreal Impact. Action from the Eastern Conference match at Orlando Citrus Bowl in Florida.
Sky Sports 3|1463949000|Football Gold|Chelsea v Tottenham Hotspur: 1993/94||0|0|Football,Soccer|Classic archive action from 1993/94 when Chelsea met Tottenham Hotspur at Stamford Bridge.(c)
Sky Sports 3|1463949900|Football Gold|Chelsea v Tottenham Hotspur: 2008 League Cup Final||0|0|Football,Soccer|Archive action from the 2008 League Cup Final, when Chelsea met Tottenham Hotspur at Wembley Stadium.(c)
Sky Sports 3|1463950500|Live MLS|Portland Timbers v Vancouver Whitecaps||0|0|Football - Club|Portland Timbers v Vancouver Whitecaps (Kick-off TBA). Coverage of the Western Conference clash at Providence Park.(c)
Sky Sports 3|1463958300|Sky Academy Sports Scholars|Sky Scholars: Jack Bateson||0|0|General Sports|A profile of the amateur boxer.(c)
Sky Sports 3|1463958900|WWE from the Vault|Big Show v Wade Barrett||0|0|Wrestling|The Big Show v Wade Barrett.(c)
Sky Sports 3|1463959800|Super Rugby Try Time|2016||0|0|Rugby League - Domestic|A round-up of all the tries, highlights and news headlines from the most recent round of the Super Rugby season.
Sky Sports 3|1463961600|Sporting Greats|Heike Drechsler||0|0|General Sports|A look at the career of former German long jumper Heike Drechsler, who is the only woman in the history of the event to win two Olympic gold medals, having triumphed in 1992 and 2000.
Sky Sports 3|1463963400|Darts Gold|WDC Finals 94/95||0|0|Darts|Highlights of the PDC World Darts Championship finals of 1994 and 1995.
Sky Sports 3|1463965200|Darts Gold|WDC Finals 96/97||0|0|Darts|Highlights of the PDC World Darts Championship finals of 1996 and 1997.
Sky Sports 3|1463967000|Time of Our Lives|Golden Arrows||0|0|General Sports|Gary Newbon talks to Phil Taylor, Mike Gregory and Tony Green about their favourite darts memories from down the years.
Sky Sports 3|1463970600|Sporting Greats|Rafael Nadal||0|0|General Sports|A profile of Rafael Nadal, who is regarded by many as the greatest clay court tennis player of all time, having won the French Open eight times. The Spaniard has been victorious in all of the other Grand Slams at least once and claimed Olympic Gold in 2008.
Sky Sports 3|1463972400|Sporting Greats|Mal Meninga||0|0|General Sports|A profile of former Australia rugby league captain Mal Meninga, a centre who was famed for his goal-kicking ability. Meninga now coaches the Queensland State of Origin team and has guided them to a record seven consecutive series victories over New South Wales.
Sky Sports 3|1463974200|Darts Gold|WDC Finals 98/99||0|0|Darts|Highlights of the PDC World Darts Championship finals of 1998 and 1999.
Sky Sports 3|1463976000|Sporting Heroes|Sporting Heroes: Peter Reid Interviews Allan Lamb||0|0|General Sports|The football manager and pundit talks to the former England cricketer about his career, which saw him as a mainstay of the Test side during the 1980s.
Sky Sports 3|1463979600|Sporting Greats|Eddy Merckx||0|0|General Sports|A look at the career of former cyclist Eddy Merckx, who won the Tour de France on five occasions, as well as recording at least two victories in each of the `five monuments', those being the Milan-San Remo, Tour of Flanders, Paris-Roubaix, Liege-Bastogne-Liege and the Giro di Lombardia.
Sky Sports 3|1463981400|Sporting Greats|Roger Federer||0|0|General Sports|A profile of Swiss tennis star Roger Federer, who has won a record 17 Grand Slam titles, including seven at Wimbledon, to cement his reputation as one of the greatest players of all time.
Sky Sports 3|1463983200|Sporting Rivalries|Argentina v Brazil||0|0|General Sports|The intense football rivalry between Argentina and Brazil, the South American nations who have won the World Cup seven times between them.
Sky Sports 3|1463985000|Sporting Rivalries|Federer v Nadal||0|0|General Sports|A look back at the epic tennis matches played between Roger Federer and Rafael Nadal.
Sky Sports 3|1463986800|Darts Gold|WDC Finals 10/11||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2010 and 2011.
Sky Sports 3|1463988600|Darts Gold|WDC Finals 02/03||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2002 and 2003.
Sky Sports 3|1463990400|Sporting Greats|Mal Meninga||0|0|General Sports|A profile of former Australia rugby league captain Mal Meninga, a centre who was famed for his goal-kicking ability. Meninga now coaches the Queensland State of Origin team and has guided them to a record seven consecutive series victories over New South Wales.
Sky Sports 3|1463992200|Sporting Greats|Lester Piggott||0|0|General Sports|A look at the career of Lester Piggott, the former jockey who had 4,493 wins, including nine Epsom Derby victories, the first of which was when he was 18 years old. Piggott initially retired at the end of the 1985 flat racing season and became a trainer, but returned as a jockey in 1990 and went on to ride for another five years.
Sky Sports 3|1463994000|Sporting Heroes|Sporting Heroes: Gary Newbon Interviews Sir Roger Bannister||0|0|General Sports|An interview with the former athlete, famous for being the first person to run a mile in under four minutes in a competitive athletics event.
Sky Sports 3|1463997600|Racing News|2016||0|0|Horse racing|Preview of race meetings across the country - including the latest betting news from today's cards.
Sky Sports 3|1463999400|Sporting Greats|Eddy Merckx||0|0|General Sports|A look at the career of former cyclist Eddy Merckx, who won the Tour de France on five occasions, as well as recording at least two victories in each of the `five monuments', those being the Milan-San Remo, Tour of Flanders, Paris-Roubaix, Liege-Bastogne-Liege and the Giro di Lombardia.
Sky Sports 3|1464001200|Super Rugby Try Time|2016||0|0|Rugby League - Domestic|A round-up of all the tries, highlights and news headlines from the most recent round of the Super Rugby season.
Sky Sports 3|1464003000|Sporting Heroes|Sporting Heroes: Greg Rutherford Interviews Lynn Davies||0|0|Athletics|The current Olympic long jump champion meets the man who won gold at the 1964 Games in Tokyo, to discuss his memories and how the sport has changed.
Sky Sports 3|1464006600|Time of Our Lives|Champion Jockeys||0|0|General Sports|Former jockeys Willie Carson, Pat Eddery and Joe Mercer look back on their careers.
Sky Sports 3|1464010200|Sporting Rivalries|USSR v USA||0|0|General Sports|A look at the basketball rivalry shared between the USSR and USA.
Sky Sports 3|1464012000|Barclays Premier League Legends|PL Legends: David Ginola||0|0|Football - Club|The Premier League career of David Ginola, the charismatic French winger who made 195 appearances during spells with Newcastle United, Tottenham Hotspur, Aston Villa and Everton.
Sky Sports 3|1464013800|Premier League Years|1997/98||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 1997/98 season, all set to a specially selected soundtrack from the time.
Sky Sports 3|1464021000|Sporting Greats|Heike Drechsler||0|0|General Sports|A look at the career of former German long jumper Heike Drechsler, who is the only woman in the history of the event to win two Olympic gold medals, having triumphed in 1992 and 2000.
Sky Sports 3|1464022800|Super Rugby Try Time|2016||0|0|Rugby League - Domestic|A round-up of all the tries, highlights and news headlines from the most recent round of the Super Rugby season.
Sky Sports 3|1464024600|Premier League 100 Club|PL 100 Club: Emile Heskey||0|0|Football - Club|The best of Emile Heskey's top-flight goals, which he scored with five different clubs - Leicester City, Liverpool, Birmingham City, Wigan Athletic and Aston Villa.
Sky Sports 3|1464026400|Cycling|The Rutland-Melton International CiCLE Classic||0|0|Cycling|The Rutland-Melton International CiCLE Classic. Action from the event that starts in Oakham and finishes in Melton Mowbray.
Sky Sports 3|1464030000|Sky Sports Boxing Gold|Anthony Joshua v Raphael Zumbano Love||0|0|Boxing|Anthony Joshua v Raphael Zumbano Love.
Sky Sports 3|1464031200|Sky Sports Boxing Gold|Anthony Joshua v Jason Gavern||0|0|Boxing|Anthony Joshua v Jason Gavern. Action from the heavyweight bout, which took place at the Metro Radio Arena in Newcastle in April 2015.
Sky Sports 3|1464032400|Sky Sports Boxing Gold|Anthony Joshua v Konstantin Airich||0|0|Boxing|Anthony Joshua v Konstantin Airich.
Sky Sports 3|1464033600|Cycling|The Rutland-Melton International CiCLE Classic||0|0|Cycling|The Rutland-Melton International CiCLE Classic. Action from the event that starts in Oakham and finishes in Melton Mowbray.
Sky Sports 3|1464037200|Premier League Years|1997/98||0|0|Football - Club|Classic games, infamous blunders and moments of skill from the 1997/98 season, all set to a specially selected soundtrack from the time.
Sky Sports 3|1464044400|Super Rugby Try Time|2016||0|0|Rugby League - Domestic|A round-up of all the tries, highlights and news headlines from the most recent round of the Super Rugby season.(n)
Sky Sports 3|1464046200|Darts Gold|WDC Finals 06/07||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2006 and 2007.(n)
Sky Sports 3|1464048000|Sporting Greats|Sergey Bubka||0|0|General Sports|A profile of Sergey Bubka, who won the gold medal at the 1988 Olympic Games in Seoul, and held the world pole vault record from 1984 to 2014.(n)
Sky Sports 3|1464049800|Sporting Greats|Michael Johnson||0|0|General Sports|A profile of Michael Johnson, the American sprinter who won four Olympic gold medals, in addition to eight golds at the World Championships. A specialist in both the 200m and 400m events, Johnson broke his own world record at the 1996 Games in Atlanta, winning the 200m final in a time of 19.32 seconds, a record which stood until the emergence of Usain Bolt.(n)
Sky Sports 3|1464051600|Sporting Greats|Heike Drechsler||0|0|General Sports|A look at the career of former German long jumper Heike Drechsler, who is the only woman in the history of the event to win two Olympic gold medals, having triumphed in 1992 and 2000.(n)
Sky Sports 3|1464053400|Sporting Greats|Usain Bolt||0|0|General Sports|A profile of Usain Bolt, the Jamaican sprinter who holds the current 100m and 200m world records and won three gold medals at the London Olympics.(n)
Sky Sports 3|1464055200|Time of Our Lives|Athletics '91||0|0|General Sports|Derek Redmond, John Regis and Kriss Akabusi look back at their gold medal-winning 4x400m relay display in the 1991 World Athletics Championships in Tokyo. Gary Newbon presents.(n)
Sky Sports 3|1464058800|Sporting Heroes|Sporting Heroes: Gary Newbon Interviews Jackie Joyner-Kersee||0|0|Athletics|The presenter talks to the former athlete about her life and career, which saw her pick up three Olympic gold medals in the heptathlon and the long jump between 1988 and 1992. She is also a four-time world champion, having topped the podium in the same events on two occasions apiece.(n)
Sky Sports 3|1464062400|Darts Gold|WDC Finals 10/11||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2010 and 2011.(n)
Sky Sports 3|1464064200|Darts Gold|WDC Finals 12/13||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2012 and 2013.(n)
Sky Sports 3|1464066000|Sporting Greats|Usain Bolt||0|0|General Sports|A profile of Usain Bolt, the Jamaican sprinter who holds the current 100m and 200m world records and won three gold medals at the London Olympics.(n)
Sky Sports 3|1464067800|Sporting Greats|Muhammad Ali||0|0|General Sports|A look back at the career of charismatic former boxer Muhammad Ali, who won the world heavyweight title on three occasions and is regarded as one of the greatest fighters of all time.(n)
Sky Sports 3|1464069600|Sporting Rivalries|Federer v Nadal||0|0|General Sports|A look back at the epic tennis matches played between Roger Federer and Rafael Nadal.(n)
Sky Sports 3|1464071400|Sporting Rivalries|Muhammad Ali v Joe Frazier||0|0|General Sports|A look at the memorable rivalry between Muhammad Ali and Joe Frazier, who fought each other on three occasions, culminating with the `Thrilla in Manila' in 1975.(n)
Sky Sports 3|1464073200|Sporting Heroes|Sporting Heroes: Denise Lewis Interviews Mary Peters||0|0|General Sports|The former heptathlete, who claimed gold in the 2000 Sydney Olympics, talks to the 1972 Olympic gold medallist, who triumphed in the pentathlon.(n)
Sky Sports 3|1464076800|Sporting Rivalries|Federer v Nadal||0|0|General Sports|A look back at the epic tennis matches played between Roger Federer and Rafael Nadal.(n)
Sky Sports 3|1464078600|Sporting Rivalries|Coe v Ovett||0|0|General Sports|A look back at the battles for supremacy on the track between Sebastian Coe and Steve Ovett.(n)
Sky Sports 3|1464080400|Cycling|The Rutland-Melton International CiCLE Classic||0|0|Cycling|The Rutland-Melton International CiCLE Classic. Action from the event that starts in Oakham and finishes in Melton Mowbray.(n)
Sky Sports 3|1464084000|Racing News|2016||0|0|Horse racing|Preview of race meetings across the country - including the latest betting news from today's cards.(n)
Sky Sports 3|1464085800|Darts Gold|WDC Finals 14/15||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2014 and 2015.(n)
Sky Sports 3|1464087600|First Utility Super League Highlights|Magic Weekend Highlights: Salford Red Devils v Widnes Vikings||0|0|Rugby League - Domestic|Salford Red Devils v Widnes Vikings. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464088500|First Utility Super League Highlights|Magic Weekend Highlights: Warrington Wolves v Castleford Tigers||0|0|Rugby League - Domestic|Warrington Wolves v Castleford Tigers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464089400|First Utility Super League Highlights|Magic Weekend Highlights: Leeds Rhinos v Wigan Warriors||0|0|Rugby League - Domestic|Leeds Rhinos v Wigan Warriors. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464090300|First Utility Super League Highlights|Magic Weekend Highlights: Wakefield Trinity Wildcats v Catalan Dragons||0|0|Rugby League - Domestic|Wakefield Trinity Wildcats v Catalan Dragons. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464091200|First Utility Super League Highlights|Magic Weekend Highlights: St Helens v Huddersfield Giants||0|0|Rugby League - Domestic|St Helens v Huddersfield Giants. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464092100|First Utility Super League Highlights|Magic Weekend Highlights: Hull FC v Hull Kingston Rovers||0|0|Rugby League - Domestic|Hull FC v Hull Kingston Rovers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464093000|Cycling|The Rutland-Melton International CiCLE Classic||0|0|Cycling|The Rutland-Melton International CiCLE Classic. Action from the event that starts in Oakham and finishes in Melton Mowbray.(n)
Sky Sports 3|1464096600|Sporting Rivalries|Romania v USSR||0|0|General Sports|A look at the gymnastics rivalry shared between Romania and USSR.(n)
Sky Sports 3|1464098400|Sky Sports Boxing Gold|Michael Gomez v Alex Arthur||0|0|Boxing|Alex Arthur v Michael Gomez. Action from the British Super-Featherweight title bout at the Meadowbank Leisure Centre in Edinburgh.(n)
Sky Sports 3|1464100200|Sky Sports Boxing Gold|Floyd Mayweather Jr v Ricky Hatton||0|0|Boxing|Floyd Mayweather Jr v Ricky Hatton. Action from the WBC Welterweight title bout at the MGM Grand in Las Vegas, which took place in 2007.(n)
Sky Sports 3|1464102000|First Utility Super League Highlights|Magic Weekend Highlights: Salford Red Devils v Widnes Vikings||0|0|Rugby League - Domestic|Salford Red Devils v Widnes Vikings. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464102900|First Utility Super League Highlights|Magic Weekend Highlights: Warrington Wolves v Castleford Tigers||0|0|Rugby League - Domestic|Warrington Wolves v Castleford Tigers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464103800|First Utility Super League Highlights|Magic Weekend Highlights: Leeds Rhinos v Wigan Warriors||0|0|Rugby League - Domestic|Leeds Rhinos v Wigan Warriors. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464104700|First Utility Super League Highlights|Magic Weekend Highlights: Wakefield Trinity Wildcats v Catalan Dragons||0|0|Rugby League - Domestic|Wakefield Trinity Wildcats v Catalan Dragons. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464105600|First Utility Super League Highlights|Magic Weekend Highlights: St Helens v Huddersfield Giants||0|0|Rugby League - Domestic|St Helens v Huddersfield Giants. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464106500|First Utility Super League Highlights|Magic Weekend Highlights: Hull FC v Hull Kingston Rovers||0|0|Rugby League - Domestic|Hull FC v Hull Kingston Rovers. Action from the Super League match at St James' Park in Newcastle.(n)
Sky Sports 3|1464107400|Cycling|The Rutland-Melton International CiCLE Classic||0|0|Cycling|The Rutland-Melton International CiCLE Classic. Action from the event that starts in Oakham and finishes in Melton Mowbray.(n)
Sky Sports 3|1464111000|Sportswomen|2016||0|0|General Sports|The biggest talking-points in the world of women's sport, including interviews and features.(n)
Sky Sports 3|1464112800|Football Gold|Liverpool v Chelsea: 2013/14||0|0|Football,Soccer|Liverpool v Chelsea from the 2013/14 season.(n)
Sky Sports 3|1464113700|Football Gold|Sunderland v Manchester United: 2013/14||0|0|Football,Soccer|Sunderland v Manchester United from the 2013/14 Premier League season.(n)
Sky Sports 3|1464114600|Football Gold|Manchester City v Manchester United: 2013/14||0|0|Football,Soccer|Manchester City v Manchester United from the 2013/14 Premier League season, which finished 4-1.(n)
Sky Sports 3|1464115500|Football Gold|Sunderland v Liverpool: 2013/14||0|0|Football,Soccer|Sunderland v Liverpool from the 2013/14 season.(n)
Sky Sports 3|1464116400|Sky Sports Boxing Gold|Michael Gomez v Alex Arthur||0|0|Boxing|Alex Arthur v Michael Gomez. Action from the British Super-Featherweight title bout at the Meadowbank Leisure Centre in Edinburgh.(n)
Sky Sports 3|1464118200|Sky Sports Boxing Gold|David Haye v Nikolai Valuev||0|0|Boxing|Nikolai Valuev v David Haye. Action from the WBA Heavyweight title bout in November 2009 at the Arena Nurnberger Versicherung in Nuremberg, Germany.(n)
Sky Sports 3|1464120000|Sky Sports Boxing Gold|Amir Khan v Andriy Kotelnik||0|0|Boxing|Andriy Kotelnik v Amir Khan. Action from the WBA Light Welterweight title bout, which took place at Manchester's MEN Arena in 2009.(n)
Sky Sports 3|1464121800|Sportswomen|2016||0|0|General Sports|The biggest talking-points in the world of women's sport, including interviews and features.(n)
Sky Sports 3|1464123600|Live Sky Poker|||0|0|Poker|Coverage of the Sky Poker Grudge Match, as a recreational player takes on one of Sky's team of professionals.(n)
Sky Sports 4|1463871600|Golf Special|An Evening with Rory McIlroy||0|0|Golf|A special event from the Irish Open, with guests including Sir Alex Ferguson and James Nesbitt.
Sky Sports 4|1463875200|PGA Tour Classic|1992 K-Mart Greater Greensboro Open||0|0|Golf|The 1992 K-Mart Greater Greensboro Open. Highlights from the Forest Oaks Country Club in Greensboro.
Sky Sports 4|1463878800|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Three||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day three of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1463882400|Golf Special|An Evening with Rory McIlroy||0|0|Golf|A special event from the Irish Open, with guests including Sir Alex Ferguson and James Nesbitt.
Sky Sports 4|1463886000|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Three||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day three of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1463889600|PGA Tour Classic|2001 Buick Classic||0|0|Golf|The 2001 Buick Classic. Archive action from the PGA Tour event at Westchester Country Club in New York.
Sky Sports 4|1463893200|PGA Tour Classic|2001 Bay Hill Invitational||0|0|Golf|The 2001 Bay Hill Invitational. Highlights from the tournament held at the Bay Hill Club and Lodge in Orlando, where defending champion Tiger Woods battled it out with Phil Mickelson for the title.
Sky Sports 4|1463896800|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Three||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day three of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1463900400|Golf Special|An Evening with Rory McIlroy||0|0|Golf|A special event from the Irish Open, with guests including Sir Alex Ferguson and James Nesbitt.
Sky Sports 4|1463904000|WWE: Smackdown|||0|0|Wrestling|Spectacular grappling action with the over-the-top stars of the States, profiling fighters causing a stir and following feuds as they spill out of the ring.
Sky Sports 4|1463907600|WWE: Experience|||0|0|Wrestling|Round-up of the latest from Raw and Smackdown, including interviews with some of the biggest stars in the sport.
Sky Sports 4|1463911200|Golf Special|An Evening with Rory McIlroy||0|0|Golf|A special event from the Irish Open, with guests including Sir Alex Ferguson and James Nesbitt.
Sky Sports 4|1463914800|WWE: Raw|||0|0|Wrestling|Wrestling action from the States with the over-the-top stars, featuring the likes of Randy Orton and John Cena. Presented by Michael Cole, John `Bradshaw' Layfield and Byron Saxton.
Sky Sports 4|1463918400|Live European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Coverage of the fourth and final day of the event, held this year at the K Club in Straffan, Co Kildare.(c)
Sky Sports 4|1463936400|Live PGA Tour Golf|2016 AT&T Byron Nelson: Day Four||0|0|Golf|The AT&T Byron Nelson. Coverage of the fourth and final day at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch is the defending champion.(c)
Sky Sports 4|1463954400|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1463958000|Golf Special|An Evening with Rory McIlroy||0|0|Golf|A special event from the Irish Open, with guests including Sir Alex Ferguson and James Nesbitt.
Sky Sports 4|1463961600|PGA Tour Classic|2003 MCI Heritage Classic||0|0|Golf|Highlights of the 2003 MCI Heritage Classic from the Harbour Town Golf Links on Hilton Head Island, South Carolina, where Justin Leonard entered as the defending champion.
Sky Sports 4|1463965200|The Sky Sports Years|1995||0|0|Sports Magazines|Action from 1995, the fifth year of Sky Sports coverage, featuring vintage moments from the time.
Sky Sports 4|1463968800|Sporting Greats|Usain Bolt||0|0|General Sports|A profile of Usain Bolt, the Jamaican sprinter who holds the current 100m and 200m world records and won three gold medals at the London Olympics.
Sky Sports 4|1463970600|Sporting Triumphs|Michael Atherton Batting for Two Days Against South Africa||0|0|General Sports|Former England cricket captain Michael Atherton relives his most memorable sporting moment, when he held firm against a South African bowling attack featuring Allan Donald in 1998.
Sky Sports 4|1463971500|Sporting Triumphs|Dennis Taylor Winning 1985 Snooker World Final||0|0|General Sports|Dennis Taylor relives his memorable world snooker championship win in 1985, when he overcame Steve Davis in a gripping final watched by more than 18 million TV viewers in the UK.
Sky Sports 4|1463972400|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1463976000|PGA Tour Classic|2000 SEI Pennsylvania Classic||0|0|Golf|The 2000 SEI Pennsylvania Classic. Action from the tournament staged at the Waynesborough Country Club in Paoli, Pennsylvania.
Sky Sports 4|1463979600|PGA Tour Classic|1996 Quad City Classic||0|0|Golf|A chance to look back at the 1996 Quad City Classic at the Oakwood Country Club in Coal Valley, Illinois.
Sky Sports 4|1463983200|Shell's Wonderful World of Golf|Annika Sorenstam v Dottie Pepper: 1996||0|0|Golf|A chance to relive the 1996 battle between Annika Sorenstam and Dottie Pepper on the Ocean Course at Kiawah Island in South Carolina. Sorenstam had 72 LPGA tournament wins to her name when she retired from golf in 2008, including 10 Majors.
Sky Sports 4|1463988600|PGA Tour Golf|2016 AT&T Byron Nelson: Day Four||0|0|Golf|The AT&T Byron Nelson. Highlights of the fourth and final day at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch was the defending champion.
Sky Sports 4|1464004800|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1464008400|Sporting Greats|Jack Nicklaus||0|0|General Sports|A look at the career of Jack Nicklaus, who is widely considered as the greatest golfer in the history of the game, after winning a total of 18 Majors. His first came at the 1962 US Open, while his most recent was the 1986 Masters, which saw him claim a sixth Green Jacket and become the oldest winner of that tournament.
Sky Sports 4|1464010200|Sporting Rivalries|The Ryder Cup||0|0|General Sports|The golfing rivalry between America and Europe, which comes to a head every two years at the Ryder Cup.
Sky Sports 4|1464012000|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1464015600|Shell's Wonderful World of Golf|Ernie Els v Nick Price: 1999||0|0|Golf|A chance to see what happened when Ernie Els clashed with Nick Price at Leopard Creek Country Club in Mpumalanga, South Africa, in 1999.
Sky Sports 4|1464021000|Sporting Greats|Jack Nicklaus||0|0|General Sports|A look at the career of Jack Nicklaus, who is widely considered as the greatest golfer in the history of the game, after winning a total of 18 Majors. His first came at the 1962 US Open, while his most recent was the 1986 Masters, which saw him claim a sixth Green Jacket and become the oldest winner of that tournament.
Sky Sports 4|1464022800|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1464026400|PGA Tour Golf|2016 AT&T Byron Nelson: Review||0|0|Golf|The AT&T Byron Nelson. Highlights of the recent event at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch was the defending champion.
Sky Sports 4|1464030000|Top 14 Rugby Union Highlights|2015/16||0|0|Rugby Union - Domestic|Action from the latest round of fixtures in France's top domestic competition.
Sky Sports 4|1464031800|Chronicles of a Champion Golfer|Greg Norman||0|0|Golf|A profile of Greg Norman.
Sky Sports 4|1464033600|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.
Sky Sports 4|1464037200|PGA Tour Golf|2016 AT&T Byron Nelson: Review||0|0|Golf|The AT&T Byron Nelson. Highlights of the recent event at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch was the defending champion.
Sky Sports 4|1464040800|Time of Our Lives|Athletics '91||0|0|General Sports|Derek Redmond, John Regis and Kriss Akabusi look back at their gold medal-winning 4x400m relay display in the 1991 World Athletics Championships in Tokyo. Gary Newbon presents.
Sky Sports 4|1464044400|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.(n)
Sky Sports 4|1464048000|PGA Tour Golf|2016 AT&T Byron Nelson: Review||0|0|Golf|The AT&T Byron Nelson. Highlights of the recent event at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch was the defending champion.(n)
Sky Sports 4|1464051600|PGA Tour Classic|1998 Mastercard Colonial||0|0|Golf|The best moments from the 1998 Mastercard Colonial at the Colonial Country Club in Texas.(n)
Sky Sports 4|1464055200|PGA Tour Classic|1993 Memorial Tournament||0|0|Golf|A chance to relive the finest moments from the 1993 Memorial Tournament at the Muirfield Village Golf Club in Ohio.(n)
Sky Sports 4|1464058800|Shell's Wonderful World of Golf|Annika Sorenstam v Dottie Pepper: 1996||0|0|Golf|A chance to relive the 1996 battle between Annika Sorenstam and Dottie Pepper on the Ocean Course at Kiawah Island in South Carolina. Sorenstam had 72 LPGA tournament wins to her name when she retired from golf in 2008, including 10 Majors.(n)
Sky Sports 4|1464064200|Sporting Rivalries|The Ryder Cup||0|0|General Sports|The golfing rivalry between America and Europe, which comes to a head every two years at the Ryder Cup.(n)
Sky Sports 4|1464066000|PGA Tour Classic|1988 Manufacturers Hanover Westchester Classic||0|0|Golf|A look back at the 1988 Manufacturers Hanover Westchester Classic at Westchester Country Club in New York. JC Snead went into the tournament as the defending champion.(n)
Sky Sports 4|1464069600|Shell's Wonderful World of Golf|Johnny Miller v Jack Nicklaus: 1997||0|0|Golf|A look back at the 1997 showdown between Johnny Miller and Jack Nicklaus at the Olympic Club in San Francisco, California. Nicklaus is the most successful man to have played the game with 18 Majors to his name, while Miller was one of the top players of the 1970s, winning the US Open in 1973 and the Open in 1976.(n)
Sky Sports 4|1464075000|Darts Gold|WDC Finals 04/05||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2004 and 2005.(n)
Sky Sports 4|1464076800|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.(n)
Sky Sports 4|1464080400|Shell's Wonderful World of Golf|Johnny Miller v Jack Nicklaus: 1997||0|0|Golf|A look back at the 1997 showdown between Johnny Miller and Jack Nicklaus at the Olympic Club in San Francisco, California. Nicklaus is the most successful man to have played the game with 18 Majors to his name, while Miller was one of the top players of the 1970s, winning the US Open in 1973 and the Open in 1976.(n)
Sky Sports 4|1464085800|Top 14 Rugby Union Highlights|2015/16||0|0|Rugby Union - Domestic|Action from the latest round of fixtures in France's top domestic competition.(n)
Sky Sports 4|1464087600|PGA Tour Golf|2016 AT&T Byron Nelson: Review||0|0|Golf|The AT&T Byron Nelson. Highlights of the recent event at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch was the defending champion.(n)
Sky Sports 4|1464091200|European Tour Golf|2016 Irish Open Hosted by the Rory Foundation: Day Four||0|0|Golf|The Irish Open Hosted by the Rory Foundation. Highlights of day four of the event, held this year at the K Club in Straffan, Co Kildare.(n)
Sky Sports 4|1464094800|PGA Tour Classic|1988 Manufacturers Hanover Westchester Classic||0|0|Golf|A look back at the 1988 Manufacturers Hanover Westchester Classic at Westchester Country Club in New York. JC Snead went into the tournament as the defending champion.(n)
Sky Sports 4|1464098400|Sporting Greats|Gary Player||0|0|General Sports|A look back at the career of South African golfer Gary Player, who won nine Majors during the 1960s and 1970s, and is the only non-American to win all four Major tournaments.(n)
Sky Sports 4|1464100200|PGA Tour Golf|2016 AT&T Byron Nelson: Review||0|0|Golf|The AT&T Byron Nelson. Highlights of the recent event at the TPC Four Seasons Resort in Irving, Texas, where Steven Bowditch was the defending champion.(n)
Sky Sports 4|1464103800|Shell's Wonderful World of Golf|Johnny Miller v Jack Nicklaus: 1997||0|0|Golf|A look back at the 1997 showdown between Johnny Miller and Jack Nicklaus at the Olympic Club in San Francisco, California. Nicklaus is the most successful man to have played the game with 18 Majors to his name, while Miller was one of the top players of the 1970s, winning the US Open in 1973 and the Open in 1976.(n)
Sky Sports 4|1464109200|MLS Round-Up Show|2016||0|0|Football - Club|A review of the latest round of Major League Soccer fixtures.(n)
Sky Sports 4|1464111000|Golfing World|2016||0|0|Golf|Magazine show, featuring news, highlights, features, tips and resort reviews, along with documentaries getting behind the scenes of the biggest events in the sport.(n)
Sky Sports 4|1464112800|Sporting Heroes|Sporting Heroes: Phil Tufnell Interviews Tony Adams||0|0|General Sports|The cricket pundit talks to the former England footballer about his career, which saw him as a mainstay of the Arsenal side during a golden period for the club.(n)
Sky Sports 4|1464116400|Top 14 Rugby Union Highlights|2015/16||0|0|Rugby Union - Domestic|Action from the latest round of fixtures in France's top domestic competition.(n)
Sky Sports 4|1464118200|Golfing World|2016||0|0|Golf|Magazine show, featuring news, highlights, features, tips and resort reviews, along with documentaries getting behind the scenes of the biggest events in the sport.(n)
Sky Sports 4|1464120000|Sporting Heroes|Sporting Heroes: Gary Newbon Interviews Mary Rand||0|0|General Sports|An interview with the 1964 Olympic long jump champion, who became the first-ever British female to win an Olympic gold medal in a track and field event.(n)
Sky Sports 4|1464123600|Golfing World|2016||0|0|Golf|Magazine show, featuring news, highlights, features, tips and resort reviews, along with documentaries getting behind the scenes of the biggest events in the sport.(n)
Sky Sports 4|1464125400|Sporting Greats|Gary Player||0|0|General Sports|A look back at the career of South African golfer Gary Player, who won nine Majors during the 1960s and 1970s, and is the only non-American to win all four Major tournaments.(n)
Sky Sports 4|1464127200|PGA Tour Classic|1988 Manufacturers Hanover Westchester Classic||0|0|Golf|A look back at the 1988 Manufacturers Hanover Westchester Classic at Westchester Country Club in New York. JC Snead went into the tournament as the defending champion.(n)
Sky Sports 5|1463873400|Football's Greatest Players|Thierry Henry||0|0|Football - International|A look back at the career of former Arsenal and France star Thierry Henry.
Sky Sports 5|1463875200|Football's Greatest International Teams|Brazil 1982||0|0|Football - International|A profile of the Brazil side that starred at the 1982 FIFA World Cup in Spain, which failed to lift the famous trophy, but delighted crowds with their style of play.
Sky Sports 5|1463877000|Football's Greatest International Teams|France 1984||0|0|Football - International|A profile of the France team that triumphed at the 1984 European Championships, featuring interviews with former players and some of the journalists that covered the tournament.
Sky Sports 5|1463878800|Football's Greatest Players|Steven Gerrard||0|0|Football - International|The career of former Liverpool and England captain Steven Gerrard.
Sky Sports 5|1463880600|Football's Greatest Players|Cristiano Ronaldo||0|0|Football - International|The career of Real Madrid and Portugal star Cristiano Ronaldo.
Sky Sports 5|1463882400|Football's Greatest Players|Luis Figo||0|0|Football - International|The career of Luis Figo, who played for Real Madrid and Barcelona, as well as excelling for Portugal.
Sky Sports 5|1463884200|Football's Greatest Players|Thierry Henry||0|0|Football - International|A look back at the career of former Arsenal and France star Thierry Henry.
Sky Sports 5|1463886000|Football's Greatest International Teams|Brazil 1982||0|0|Football - International|A profile of the Brazil side that starred at the 1982 FIFA World Cup in Spain, which failed to lift the famous trophy, but delighted crowds with their style of play.
Sky Sports 5|1463887800|Football's Greatest International Teams|France 1984||0|0|Football - International|A profile of the France team that triumphed at the 1984 European Championships, featuring interviews with former players and some of the journalists that covered the tournament.
Sky Sports 5|1463889600|Time of Our Lives|SW19 Ladies||0|0|General Sports|Wimbledon ladies' stars Virginia Wade, Ann Jones and Angela Mortimer reminisce about their glittering careers on the grass courts of the All England Club. Presented by Gary Newbon.
Sky Sports 5|1463893200|Indian Premier League|Gujarat Lions v Mumbai Indians||0|0|Cricket - Domestic|Gujarat Lions v Mumbai Indians. Action from the Twenty20 match, which took place at Green Park in Kanpur.
Sky Sports 5|1463909400|Darts Gold|WDC Finals 14/15||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2014 and 2015.
Sky Sports 5|1463911200|Live Indian Premier League|Kolkata Knight Riders v Sunrisers Hyderabad||0|0|Cricket - Domestic|Kolkata Knight Riders v Sunrisers Hyderabad. All the action from Eden Gardens, where the lucrative Twenty20 competition continues.
Sky Sports 5|1463925600|Live Indian Premier League|Delhi Daredevils v Royal Challengers Bangalore||0|0|Cricket - Domestic|Delhi Daredevils v Royal Challengers Bangalore. Coverage of the group-stage match in the Twenty20 competition, from Feroz Shah Kotla.
Sky Sports 5|1463941800|Football's Greatest Players|Clarence Seedorf||0|0|Football - International|The career of former AC Milan and Netherlands star Clarence Seedorf.
Sky Sports 5|1463943600|WWE Special|The John Cena Experience||0|0|Wrestling|An insight into the life of John Cena, who has claimed the WWE Championship on 10 occasions and won 19 titles in total, featuring a look at his preparations for wrestling bouts and his life away from the sport.
Sky Sports 5|1463947200|WWE: Late Night - Raw|||0|0|Wrestling|Wrestling action from the States with the over-the-top stars, featuring the likes of Randy Orton and John Cena. Presented by Michael Cole.
Sky Sports 5|1463950800|WWE: Late Night - Smackdown|||0|0|Wrestling|Spectacular wrestling action with the over-the-top stars of the States, profiling fighters causing a stir and following feuds as they spill out of the ring.
Sky Sports 5|1463954400|WWE Main Event|||0|0|Wrestling|Michael Cole and Byron Saxton present wrestling action featuring stars from the WWE roster.
Sky Sports 5|1463958000|Football's Greatest Players|Alan Shearer||0|0|Football - International|The career of former Newcastle United and England striker Alan Shearer.
Sky Sports 5|1463959800|Football's Greatest Players|Lionel Messi||0|0|Football - International|The career of Barcelona and Argentina star Lionel Messi.
Sky Sports 5|1463961600|Football's Greatest Players|Andres Iniesta||0|0|Football - International|The career of Barcelona and Spain star Andres Iniesta, who has been one of the leading players in the world over the past decade.
Sky Sports 5|1463963400|Football's Greatest Players|Ryan Giggs||0|0|Football - International|The career of former Manchester United and Wales star Ryan Giggs, who is the most decorated player in English football history.
Sky Sports 5|1463965200|Time of Our Lives|Wigan Warriors||0|0|General Sports|Former Wigan Warriors stars Shaun Edwards, Ellery Hanley and Martin Offiah look back on their time with the club. Gary Newbon presents.
Sky Sports 5|1463968800|Football's Greatest Teams|Nottingham Forest||1|13|Football,Soccer|A look at Brian Clough's Nottingham Forest side from the mid to late 1970s, featuring archive footage and interviews with Peter Shilton and Martin O'Neill.
Sky Sports 5|1463970600|Football's Greatest Teams|Santos||0|0|Football,Soccer|A look at the Santos side of the 1960s, which included the likes of Zito, Carlos Alberto and Pele.
Sky Sports 5|1463972400|Football's Greatest Teams|Red Star Belgrade||0|0|Football,Soccer|A look at 1991 European Cup-winning Red Star Belgrade side, which included such stars as Darko Pancev, Robert Prosinecki and Sinisa Mihajlovic.
Sky Sports 5|1463974200|Football's Greatest Teams|Liverpool||1|11|Football,Soccer|A look at the success enjoyed by Liverpool during the 1970s and 80s, featuring interviews with the likes of Kenny Dalglish, Alan Hansen and Graeme Souness.
Sky Sports 5|1463976000|Time of Our Lives|Grapple Greats||0|0|General Sports|Gary Newbon talks to former British wrestlers, including Banger Walsh, Mark `Rollerball' Rocco and Mick McManus.
Sky Sports 5|1463979600|Good Morning Sports Fans|||0|0|General Sports|News and views on today's early stories, a look at the back pages, a tip on today's racing and a sporting weather forecast.
Sky Sports 5|1463983200|Good Morning Sports Fans|||0|0|General Sports|News and views on today's early stories, a look at the back pages, a tip on today's racing and a sporting weather forecast.
Sky Sports 5|1463986800|Good Morning Sports Fans|||0|0|General Sports|News and views on today's early stories, a look at the back pages, a tip on today's racing and a sporting weather forecast.
Sky Sports 5|1463990400|Time of Our Lives|Speedway Stars||0|0|General Sports|Michael Lee, Gary Havelock and Mark Loram reminisce about their speedway careers. Presented by Gary Newbon.
Sky Sports 5|1463994000|Super Rugby Try Time|2016||0|0|Rugby League - Domestic|A round-up of all the tries, highlights and news headlines from the most recent round of the Super Rugby season.
Sky Sports 5|1463995800|Football's Greatest Players|Dennis Bergkamp||0|0|Football - International|The career of former Arsenal and Netherlands star Dennis Bergkamp.
Sky Sports 5|1463997600|Time of Our Lives|Olympics 1964||0|0|General Sports|Former athletes Lynn Davies, Ken Matthews and Ann Packer reminisce about their performances at the 1964 Tokyo Olympics, which saw them win gold medals in the men's long jump, men's 20km walk and the women's 800m respectively.
Sky Sports 5|1464001200|Football's Greatest Players|Marco van Basten||0|0|Football - International|The career of former Ajax and Netherlands star Marco van Basten, who went on to manage his country after retiring as a player. The prolific striker boasted an outstanding scoring record, and will be best remembered for his wonder goal in the final of the 1988 European Championships.
Sky Sports 5|1464003000|Football's Greatest Players|Paolo Maldini||0|0|Football - International|The career of former AC Milan and Italy star Paolo Maldini, who spent his entire 25-year career with the Milanese club, which saw him win the European Cup on five occasions and the Serie A title seven times.
Sky Sports 5|1464004800|Major League Soccer|MLS Highlights: Portland Timbers v Vancouver Whitecaps||0|0|Football - Club|Portland Timbers v Vancouver Whitecaps. Action from the Western Conference clash at Providence Park.
Sky Sports 5|1464012000|Major League Soccer|MLS Highlights: Los Angeles Galaxy v San Jose Earthquakes||0|0|Football - Club|Los Angeles Galaxy v San Jose Earthquakes. Action from the Western Conference clash at StubHub Centre.
Sky Sports 5|1464019200|WWE: Raw|||0|0|Wrestling|Wrestling action from the States with the over-the-top stars, featuring the likes of Randy Orton and John Cena. Presented by Michael Cole, John `Bradshaw' Layfield and Byron Saxton.
Sky Sports 5|1464026400|Football's Greatest Managers|Fabio Capello||0|0|Football,Soccer|A profile of former England manager Fabio Capello, whose managerial career has also seen him at the helm of some of European football's top clubs, including AC Milan, Real Madrid, AS Roma and Juventus. Capello also had a distinguished playing career that saw him win 32 caps for his country.
Sky Sports 5|1464028200|Fantasy Football Club - The Highlights|2015/16||0|0|Football - Club|Max Rushden and Paul Merson look back on highlights of the show, which focusses on key fantasy football issues, and features studio guests.
Sky Sports 5|1464030000|Sporting Heroes|Sporting Heroes: Ravi Bopara Interviews Sol Campbell||0|0|Football,Soccer|The England all-rounder speaks to the former Arsenal and Tottenham Hotspur defender, who was part of the Gunners' `Invincibles' of 2003/04 and also played 73 times for England.
Sky Sports 5|1464033600|Football's Greatest Players|Ryan Giggs||0|0|Football - International|The career of former Manchester United and Wales star Ryan Giggs, who is the most decorated player in English football history.
Sky Sports 5|1464035400|Fantasy Football Club - The Highlights|2015/16||0|0|Football - Club|Max Rushden and Paul Merson look back on highlights of the show, which focusses on key fantasy football issues, and features studio guests.
Sky Sports 5|1464037200|WWE: Late Night - Raw|||0|0|Wrestling|Wrestling action from the States with the over-the-top stars, featuring the likes of Randy Orton and John Cena. Presented by Michael Cole.
Sky Sports 5|1464040800|Sporting Heroes|Sporting Heroes: Gary Newbon Interviews Jackie Joyner-Kersee||0|0|Athletics|The presenter talks to the former athlete about her life and career, which saw her pick up three Olympic gold medals in the heptathlon and the long jump between 1988 and 1992. She is also a four-time world champion, having topped the podium in the same events on two occasions apiece.
Sky Sports 5|1464044400|Darts Gold|WDC Finals 04/05||0|0|Darts|Highlights of the PDC World Darts Championship finals of 2004 and 2005.(n)
Sky Sports 5|1464046200|Football's Greatest Managers|Fabio Capello||0|0|Football,Soccer|A profile of former England manager Fabio Capello, whose managerial career has also seen him at the helm of some of European football's top clubs, including AC Milan, Real Madrid, AS Roma and Juventus. Capello also had a distinguished playing career that saw him win 32 caps for his country.(n)
Sky Sports 5|1464048000|Live WWE: Late Night - Raw|||0|0|Wrestling|Wrestling coverage from the States with the over-the-top stars, featuring the likes of Randy Orton and John Cena. Presented by Michael Cole.(n)
Sky Sports 5|1464059700|WWE from the Vault|Rey Mysterio and Alex Riley v The Miz and Jack Swagger||0|0|Wrestling|Rey Mysterio and Alex Riley v The Miz and Jack Swagger. Action from the tag team bout which took place in June 2011.(n)
Sky Sports 5|1464060600|WWE from the Vault|Alberto Del Rio v R Truth v Rey Mysterio||0|0|Wrestling|Alberto Del Rio v R Truth v Rey Mysterio. A chance to relive the triple threat match staged on an episode of Raw in July 2011. The contest was used to determine the number one contender to battle for the WWE Championship at Money in the Bank.(n)
Sky Sports 5|1464061500|WWE from the Vault|Rey Mysterio v The Miz||0|0|Wrestling|Rey Mysterio v the Miz. Action from the bout that took place in July 2011.(n)
Sky Sports 5|1464062400|Football's Greatest Teams|Benfica||1|8|Football,Soccer|A look at the success achieved by Benfica during the 1960s, featuring archive footage and interviews with the likes of Eusebio and Antonio Simoes.(n)
Sky Sports 5|1464064200|Football's Greatest Teams|Ajax||1|7|Football,Soccer|A look at the successful Ajax team of the early 1970s, featuring interviews with the likes of Rinus Michels, Johan Cruyff and Sjaak Swart.(n)
Sky Sports 5|1464066000|Good Morning Sports Fans|||0|0|General Sports|News and views on today's early stories, a look at the back pages, a tip on today's racing and a sporting weather forecast.(n)
Sky Sports 5|1464069600|Good Morning Sports Fans|||0|0|General Sports|News and views on today's early stories, a look at the back pages, a tip on today's racing and a sporting weather forecast.(n)
Sky Sports 5|1464073200|Good Morning Sports Fans|||0|0|General Sports|News and views on today's early stories, a look at the back pages, a tip on today's racing and a sporting weather forecast.(n)
Sky Sports 5|1464076800|Time of Our Lives|The Middleweights||0|0|General Sports|Three British former middleweight boxers, Alan Minter, Herol `Bomber' Graham and Tony Sibson, reminisce about their careers. Minter held two versions of the world title before losing to `Marvellous' Marvin Hagler at Wembley Arena, Graham had three unsuccessful challenges for world honours, as did Sibson, one of which was against Hagler.(n)
Sky Sports 5|1464080400|Football's Greatest Players|Steven Gerrard||0|0|Football - International|The career of former Liverpool and England captain Steven Gerrard.(n)
Sky Sports 5|1464082200|Football's Greatest Players|Cristiano Ronaldo||0|0|Football - International|The career of Real Madrid and Portugal star Cristiano Ronaldo.(n)
Sky Sports 5|1464084000|Time of Our Lives|Olympics Mexico City 1968||0|0|General Sports|British competitors David Hemery, Sheila Sherwood and David Broome reminisce about their performances at the 1968 Mexico City Olympics. Hemery won gold in the 400m hurdles, while Sherwood claimed a silver in the long jump, and Broome finished third in the individual show jumping discipline.(n)
Sky Sports 5|1464087600|Sporting Heroes|Sporting Heroes: Dickie Davies Interviews Tom Finney||0|0|General Sports|A chat with the former football player, who played for Preston North End in the 1940s, 50s and 60s, and represented England on 76 occasions.(n)
Sky Sports 5|1464091200|Sporting Heroes|Sporting Heroes: Bob Wilson Interviews Gordon Banks||0|0|General Sports|The former Arsenal goalkeeper interviews the man who played in goal for England in the 1966 World Cup, and became infamous for his save four years later against Brazil.(n)
Sky Sports 5|1464094800|Time of Our Lives|The Featherweights||0|0|General Sports|Former featherweight boxers Barry McGuigan, Colin McMillan and Steve Robinson reminisce about their careers, which saw all three of them earn world titles.(n)
Sky Sports 5|1464098400|Football's Greatest Players|Ferenc Puskas||0|0|Football - International|The career of former Real Madrid and Hungary star Ferenc Puskas, who is regarded as one of the finest goalscorers in the history of the sport, and an integral part of the 'Magnificent Magyars' team of the 1950s that became the first overseas team to beat England at Wembley Stadium.(n)
Sky Sports 5|1464100200|Football's Greatest Players|George Best||0|0|Football - International|The life and career of the former Manchester United and Northern Ireland star George Best, who won the European Cup and was named European player of the year during his time with the Red Devils.(n)
Sky Sports 5|1464102000|Football's Greatest Players|Diego Maradona||0|0|Football - International|The career of former Napoli and Argentina star Diego Maradona, who is widely considered by football fans around the world as a rival to Pele for the accolade of greatest ever player.(n)
Sky Sports 5|1464103800|Football's Greatest Players|Pele||0|0|Football - International|The career of former Santos and Brazil star Pele, who is regarded by many as the greatest player of all time. After breaking into the Santos first team at 15 years of age, he made his first appearance for the national side just one year later and helped his country succeed at the 1958 World Cup in Sweden aged 17.(n)
Sky Sports 5|1464105600|WWE: Smackdown|||0|0|Wrestling|Spectacular grappling action with the over-the-top stars of the States, profiling fighters causing a stir and following feuds as they spill out of the ring.(n)
Sky Sports 5|1464112800|Football's Greatest Managers|Rinus Michels||0|0|Football,Soccer|A profile of former Ajax, Netherlands and Barcelona manager Rinus Michels, who was widely credited with the invention of `Total Football' and whose major honours included the European Championship, the European Cup, four Dutch titles and one La Liga.(n)
Sky Sports 5|1464114600|Fantasy Football Club - The Highlights|2015/16||0|0|Football - Club|Max Rushden and Paul Merson look back on highlights of the show, which focusses on key fantasy football issues, and features studio guests.(n)
Sky Sports 5|1464116400|MLS Round-Up Show|2016||0|0|Football - Club|A review of the latest round of Major League Soccer fixtures.(n)
Sky Sports 5|1464118200|Jamie Vardy: Record Breaker|||0|0|Football - Club|A look back at the Leicester City striker's recent goalscoring achievement from earlier in the season, which saw him find the back of the net in 11 consecutive Premier League games.(n)
Sky Sports 5|1464120000|Fantasy Football Club - The Highlights|2015/16||0|0|Football - Club|Max Rushden and Paul Merson look back on highlights of the show, which focusses on key fantasy football issues, and features studio guests.(n)
Sky Sports 5|1464121800|City Slickers|||0|0|General Sports|Geoff Shreeves presents a look at the rise of Manchester City since they were bought by the Abu Dhabi United Group for Development and Investment.(n)
Sky Sports 5|1464123600|WWE: Late Night - Smackdown|||0|0|Wrestling|Spectacular wrestling action with the over-the-top stars of the States, profiling fighters causing a stir and following feuds as they spill out of the ring.(n)
Sky Sports 5|1464127200|Football's Greatest Managers|Rinus Michels||0|0|Football,Soccer|A profile of former Ajax, Netherlands and Barcelona manager Rinus Michels, who was widely credited with the invention of `Total Football' and whose major honours included the European Championship, the European Cup, four Dutch titles and one La Liga.(n)
Sky Sports 5|1464129000|Football's Greatest Managers|Mario Zagallo||0|0|Football,Soccer|A profile of Mario Zagallo, who won the World Cup as a player in 1958 and 1962, as a manager in 1970 and as an assistant coach in 1994, making him the only man to have achieved all three feats.(n)
Sky Sports F1|1463874300|Architects of F1|Flavio Briatore||0|0|Formula One|A profile of Flavio Briatore.
Sky Sports F1|1463877900|Tales from the Vault|Story of 1984||0|0|Formula One|A look back at the 1984 season.
Sky Sports F1|1463881500|Inside Mercedes|||0|0|Formula One|A look at the reigning constructors' world champions.
Sky Sports F1|1463882400|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463886000|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463889600|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463893200|Legends of F1|Legends of F1 - Mika Hakkinen||0|0|Formula One|A profile of Finnish driver Mika Hakkinen, who became world champion in 1998 and successfully defended his title the following year.
Sky Sports F1|1463896800|Legends of F1|Legends of F1 - John Surtees||0|0|Formula One|Steve Rider interviews John Surtees, the only man to have won world championships on two and four wheels.
Sky Sports F1|1463900400|F1 Midweek Report|2016 Spanish Grand Prix: Review||0|0|Formula One|A review of the Spanish Grand Prix.
Sky Sports F1|1463902200|Formula 1|2016 Australian Grand Prix: Standalone Race||0|0|Formula One|The Australian Grand Prix. A chance to see the opening round of the season at Albert Park, Melbourne, as Lewis Hamilton began his defence of the title.
Sky Sports F1|1463910300|Ted's Notebook|2016 Australia: Race||0|0|Formula One|Ted Kravitz offers his thoughts on the Australian Grand Prix.
Sky Sports F1|1463911200|Formula 1|Bahrain Grand Prix 2016: Standalone Race||0|0|Formula One|The Bahrain Grand Prix. A chance to see the second round of the season at the Bahrain International Circuit in Sakhir.
Sky Sports F1|1463919300|Ted's Notebook|2016 Bahrain: Race||0|0|Formula One|Ted Kravitz offers his thoughts on the race from Bahrain.
Sky Sports F1|1463920200|Formula 1|2016 Chinese Grand Prix: Standalone Race||0|0|Formula One|The Chinese Grand Prix. Another chance to see the third round of the season at the Shanghai International Circuit.
Sky Sports F1|1463928300|Ted's Notebook|2016 China: Race||0|0|Formula One|Ted Kravitz offers his thoughts on the Chinese Grand Prix.
Sky Sports F1|1463929200|Formula 1|2016 Russian Grand Prix: Standalone Race||0|0|Formula One|The Russian Grand Prix. A chance to see the fourth round of the season at the Sochi Autodrom.
Sky Sports F1|1463937300|Ted's Notebook|2016 Russian Grand Prix: Race||0|0|Formula One|Ted Kravitz offers his thoughts on the Russian Grand Prix.
Sky Sports F1|1463938200|Formula 1|2016 Spanish Grand Prix: Standalone Race||0|0|Formula One|The Spanish Grand Prix. A chance to see the fifth round of the season at the Circuit de Catalunya in Barcelona, where Nico Rosberg was victorious last year.
Sky Sports F1|1463946300|Ted's Notebook|2016 Spain: Race||0|0|Formula One|Ted Kravitz offers his thoughts on the Spanish Grand Prix.
Sky Sports F1|1463947200|F1 Classic Races|1992 Monaco Grand Prix||0|0|Formula One|The 1992 Monaco Grand Prix.
Sky Sports F1|1463949900|F1 Classic Races|1993 Monaco Grand Prix||0|0|Formula One|The 1993 Monaco Grand Prix.
Sky Sports F1|1463952600|F1 Midweek Report|2016 Spanish Grand Prix: Review||0|0|Formula One|A review of the Spanish Grand Prix.
Sky Sports F1|1463954400|Tales from the Vault|Family Dynasties||0|0|Formula One|A look at family dynasties, featuring the likes of Michael and Ralf Schumacher, Graham and Damon Hill, and Gilles and Jacques Villeneuve.
Sky Sports F1|1463958000|Architects of F1|Flavio Briatore||0|0|Formula One|A profile of Flavio Briatore.
Sky Sports F1|1463961600|Legends of F1|Legends of F1 - Frank Williams||0|0|Formula One|A profile of Frank Williams, the founder and team principal of the Williams F1 Formula One racing team.
Sky Sports F1|1463965200|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463968800|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463972400|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463976000|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463979600|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463983200|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463986800|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463990400|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463994000|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1463997600|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1464001200|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1464004800|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1464008400|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.
Sky Sports F1|1464011100|Formula 1|2016 Chinese Grand Prix: Standalone Race||0|0|Formula One|The Chinese Grand Prix. Another chance to see the third round of the season at the Shanghai International Circuit.
Sky Sports F1|1464019200|Legends of F1|Legends of F1 - Niki Lauda||0|0|Formula One|An interview with three-time world champion Niki Lauda.
Sky Sports F1|1464022800|Legends of F1|Legends of F1 - Mika Hakkinen||0|0|Formula One|A profile of Finnish driver Mika Hakkinen, who became world champion in 1998 and successfully defended his title the following year.
Sky Sports F1|1464026400|Tales from the Vault|Teammates||0|0|Formula One|Steve Rider is joined by Christian Horner and Nigel Mansell to discuss the biggest rivalries between F1 team-mates.
Sky Sports F1|1464030000|Tales from the Vault|Underdogs||0|0|Formula One|A look at underdogs who have succeeded in Formula One, including Damon Hill, John Watson and Pat Symonds.
Sky Sports F1|1464033600|F1 Classic Races|2003 Monaco Grand Prix||0|0|Formula One|The 2003 Monaco Grand Prix.
Sky Sports F1|1464041700|Formula 1|2016 Spanish Grand Prix: Highlights||0|0|Formula One|The Spanish Grand Prix. Action from the fifth round of the season at the Circuit de Catalunya in Barcelona.
Sky Sports F1|1464045300|Ted's Notebook|2016 Spain: Race||0|0|Formula One|Ted Kravitz offers his thoughts on the Spanish Grand Prix.(n)
Sky Sports F1|1464046200|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464048000|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464051600|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464055200|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464058800|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464062400|The Home of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464066000|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464069600|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464073200|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464076800|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464080400|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464084000|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464087600|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464091200|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464094800|The Home Of Formula One|||0|0|Formula One|The lowdown on Sky's coverage of the Formula One season.(n)
Sky Sports F1|1464097500|Formula 1|2016 Russian Grand Prix: Standalone Race||0|0|Formula One|The Russian Grand Prix. A chance to see the fourth round of the season at the Sochi Autodrom.(n)
Sky Sports F1|1464105600|F1 Midweek Report|2016 Spanish Grand Prix: Review||0|0|Formula One|A review of the Spanish Grand Prix.(n)
Sky Sports F1|1464107400|Architects of F1|Gordon Murray||0|0|Formula One|A profile of Gordon Murray.(n)
Sky Sports F1|1464111000|Formula 1|Australian F1 GP Best Bits: 2016||0|0|Formula One|A chance to relive some of the best moments from the Australian Grand Prix.(n)
Sky Sports F1|1464112800|Formula 1|Bahrain F1 GP Best Bits: 2016||0|0|Formula One|A chance to relive some of the best moments from the Bahrain Grand Prix.(n)
Sky Sports F1|1464114600|Formula 1|Chinese F1 GP Best Bits: 2016||0|0|Formula One|A chance to relive some of the best moments from the Chinese Grand Prix.(n)
Sky Sports F1|1464116400|Formula 1|Russian F1 GP Best Bits: 2016||0|0|Formula One|A look back at the key moments from the Russian Grand Prix.(n)
Sky Sports F1|1464118200|Formula 1|Spanish F1 GP Best Bits: 2016||0|0|Formula One|A chance to relive some of the best moments from the Spanish Grand Prix.(n)
Sky Sports F1|1464120000|F1 Classic Races|2008 Monaco Grand Prix||0|0|Formula One|The 2008 Monaco Grand Prix.(n)
Sky Sports F1|1464129000|Architects of F1|Jo Ramirez||0|0|Formula One|A profile of Jo Ramirez.(n)
DR1|1463868000|Amerikansk komediedrama fra 1987||1987|0|0||<h2 class='program-small-desc'>Amerikansk komediedrama fra 1987Amerikansk komediedrama fra 1987.Politimanden Burt Simpson erfarer, at han kun har kort tid tilbage at leve i. Burt beslutter sig for at blive dræbt på jobbet, så hans familie kan få udbetalt hans livsforsikring. Pludselig har stationen fået sig en ny superstrømer, der frygtløst kaster sig ud i de mest vanvittige situationer. Burt Simpson: Dabney Coleman. Ernie Dills: Matt Frewer. Carolyn: Teri Garr. Instruktion: Gregg Champion. Genre : Film. Year : 1987(n)
DR1|1463868900|Engelsk erotisk komedie fra 1994||1994|0|0||<h2 class='program-small-desc'>Engelsk erotisk komedie fra 1994Engelsk erotisk komedie fra 1994.Præsten Anthony Campion og hans kone Estella kommer på besøg hos den frisindede maler Norman Lindsay. Mens præsten forsøger at få Norman til at modere et forargeligt billede, tilbringer Estella tiden med malerens tre fordomsfri modeller. I starten forarges hun over de evigt nøgne piger, men sådan fortsætter det ikke. Anthony Campion: Hugh Grant. Estella Campion: Tara Fitzgerald. Norman Lindsay: Sam Neill. Sheela: Elle MacPherson. Instruktion: John Duigan. (t). Genre : Film. Year : 1993
DR1|1463874300|Amerikansk katastrofefilm fra 2009||2009|0|0||<h2 class='program-small-desc'>Amerikansk katastrofefilm fra 2009Amerikansk katastrofefilm fra 2009.Et voldsomt jordskælv har lavet en revne i Jordens skorpe. En revne, der bliver gradvist større. Seismologen Amy Lee og minøren Charley Baxter kommer på noget af en opgave, da de bliver sat til at finde ud af, hvilken vej revnen bevæger sig og at advare befolkningen, før det er for sent. Amy Lee: Brittany Murphy. Charley Baxter: Eriq La Salle. Dan Lane: Justin Hartley. Instruktion: David Michael Latt. (t). Genre : Film. Year : 2011
DR1|1463879400|Amerikansk komediedrama fra 1987||1987|0|0||<h2 class='program-small-desc'>Amerikansk komediedrama fra 1987Amerikansk komediedrama fra 1987.Politimanden Burt Simpson erfarer, at han kun har kort tid tilbage at leve i. Burt beslutter sig for at blive dræbt på jobbet, så hans familie kan få udbetalt hans livsforsikring. Pludselig har stationen fået sig en ny superstrømer, der frygtløst kaster sig ud i de mest vanvittige situationer. Burt Simpson: Dabney Coleman. Ernie Dills: Matt Frewer. Carolyn: Teri Garr. Instruktion: Gregg Champion. (t). Genre : Film. Year : 1987
DR1|1463884800|Udsendelsesophør|||0|0||Udsendelsesophør
DR1|1463890200|Dyst i haven (4:8)||2014|0|0||Der er syv deltagere tilbage! Sveriges største haveentusiaster er i gang med en sand kamp - mod ukrudt, mod forskellige uønskede smådyr, mod plantesygdomme og meget andet - men først og fremmest skal de i kamp mod hinanden, for hvem er den allerbedste, hvem skaber den smukkeste og mest spændende have, kort sagt: hvem er "Mesteren". Juryen består af tre meget kompetente dommere med hver deres speciale, og alt kommer til at foregå i skarp, men venskabelig konkurrence. De, der klarer dommernes opgaver bedst, går videre - men i hvert afsnit er der en, der må forlade det hyggelige selskab. Nordvision fra Sverige. (t). Episode : 4:8. Genre : Underholdning. Year : 2014
DR1|1463893800|Dyrebørnenes første tid (1:5)||2012|0|0||Naturserie fra BBC fra 2012.I maj dukker en brun bjørn op fra vinterhiet sammen med tre bittesmå unger, der for første gang kigger på verden omkring sig. Fra nu af vil deres liv dreje sig om to ting: at beskytte sig selv mod fare og en konstant kamp for at finde føde. De dybe skove er fulde af udfordringer som rovdyr, elementernes rasen og ikke mindst mennesker. De tre bjørneunger følger i hælene på deres mor og må være utrolig lærenemme for at kunne overleve det barske liv i vildmarken i den første måned af deres liv, hvor de er allermest sårbare. (t). Episode : 1:5. Genre : Dokumentar. Year : 2012
DR1|1463896800|Kæmpe havaborren||2013|0|0||Japansk naturprogram fra 2013. (t). Genre : Dokumentar. Year : 2013
DR1|1463899800|Verdens vildeste øer - Hebriderne (5:5)||2012|0|0||Hollandsk naturserie fra 2012.Verdens øer kan være hjemsted for nogle af de mest dramatiske landskaber og det mest fantastiske dyreliv. Mange tusinde års isolation har virket som brændstof på den naturlige udvælgelse, det vil sige tilpasningen til de særlige naturforhold, og har ikke alene fået de mest besynderlige væsner til at trives og overleve, men har også ført til en udvikling af nye arter specialiseret i at overleve de særlige naturforhold netop der. (t). Episode : 5:5. Genre : Natur & Miljø. Year : 2012
DR1|1463903100|Hvordan bliver man en vild elefant||2013|0|0||Canadisk naturprogram fra 2013.Den lille forældreløse elefantunge Sities har tilbragt de sidste tre år på elefantbørnehjemmet i Kenya og er ved at være gammel nok til at skulle sige farvel til børnehaven og drage syd på til den næste fase i sin tilbagevenden til naturen. I en beskyttet del af Tsavo Nationalpark følger vi Sities gennem de daglige lektioner i uafhængighed og forsigtige tilnærmelser til andre vilde elefanter. Men det tager lang tid, og det er ikke helt problemfrit! (t). Genre : Dokumentar. Year : 2013
DR1|1463905800|Spis og spar (6:6)|||0|0||Katrine og Ulrik bor i Ubby, lidt uden for Kalundborg. Ulrik er manden bag gryderne, og han elsker fløde og bacon,- og ikke grøntsager. Katrine derimod, kunne godt tænke sig at få lidt mere grønt ind i de sædvanlige retter og har også et ønske om at være lidt mere involveret i madlavningen. Men vil Ulrik give plads til Katrines ønsker og kan parret spare nok penge, til at tage hele familien med på en sommerhustur til Skagen? (t). Episode : 6:6. Genre : Fritid & Livsstil. Year : 2016
DR1|1463908500|Dronning Elizabeth - 60 år på tronen (3:3)||2012|0|0||Dokumentarserie fra BBC fra 2012.Den britiske journalist Andrew Marr, der i anledning af dronning Elizabeth den andens 60 års regeringsjubilæum har fået tilladelse til at følge dronningen gennem halvandet år, fortæller her om de afgørende øjeblikke i dronningens regeringstid, begyndende med sin tronbestigelse i 1952, og kroningen 16 måneder senere. Marr undersøger også det til tider meget anspændte forhold mellem den kongelige familie og medierne, og benytter et statsbesøg i Australien til at se på det mange mener er dronningens mest varige præstation, nemlig, at det er lykkedes dronning Elizabeth at holde sammen på Commonwealth. Og så fortæller alle de voksne børnebørn for første gang om, hvordan de opfatter deres jubilerende bedstemor. (t). Episode : 3:3. Genre : Dokumentar. Year : 2012
DR1|1463911800|Krøniken (10)||2004|0|0||- en tv-fortælling af Stig Thorsboe fra 2004.1957. Søs er netop kommet tilbage fra et besøg hos Erik i New York, da problemer på Bella gør, at belastningen bliver for meget for Kaj Holger - hele familien bliver involveret i en midlertidig løsning af den kritiske situation. Palle bliver opfordret til at stille op som folketingskandidat og må tage på besøg i Kjellerup-kredsen, som bestemt også er interesseret i den mulige kandidats kone. Der er gang i sagerne hjemme hos Børge og Karen, hvor Emma er i blomstrende pubertet, mens Ida stille og roligt forbedrer sin arbejdssituation på forlaget betydeligt. Medvirkende. Ida: Anne Louise Hassing. Erik: Ken Vedsegaard. Palle: Anders W. Berthelsen. Søs: Maibritt Saerens. Kaj Holger: Waage Sandø. Karin: Stina Ekblad. Karen: Pernille Højmark. Børge: Dick Kaysø. Vang: Finn Nielsen. Berg: John Hahn-Petersen. Sander: Thomas Mørk. Endvidere. Michael Hasselflug, Peter Hesse Overgaard, Christian Mosbæk, Anette Støvelbæk, Ole Thestrup, Bjarne Henriksen, Jacob Haugaard, Hanne Windfeld, Gladis H. Frendø, Andreas Berg Nielsen, Nis Bank-Mikkelsen, Steen Stig Lommer, Bodil Lassen, Rosa K. Frederiksen og Poul Jørgensen. Manuskript: Stig Thorsboe og Hanna Lundblad. Instruktion: Charlotte Sieling. Foto: Jørgen Johansson, dff. Scenografi: Kirsten Koch. Musik: Jacob Groth. Sendt første gang 7.3.04 (t). Episode : 10. Genre : Serier. Year : 2003. .
DR1|1463915400|UEFA EM 2016: Vejen til Frankrig|||0|0||UEFA EM 2016: Vejen til Frankrig
DR1|1463916840|OBS|||0|0||Oplysning til borgerne om samfundet. (t). Genre : Ukategoriseret. Year : 2016
DR1|1463917200|Lewis: Soning||2007|0|0||Engelsk krimi fra 2007.Rachel Mallory, mor til to og tilsyneladende lykkeligt gift, findes hængt i sit hjem. Lewis nægter at tro, at der er tale om selvmord, så han beslutter sig for at efterforske sagen som en mordsag - stik mod alle ordrer. Et meget usædvanligt forhold mellem to vennepar viser sig at være nøglen til gådens løsning. Lewis: Kevin Whately. Hathaway: Laurence Fox. Hugh Mallory: James Wilby. Instruktion: Dan Reed. (t). Genre : Serier. Year : 2006
DR1|1463922900|Hercule Poirot: Hollow-mysteriet||2003|0|0||Engelsk krimi fra 2003.Poirot er fascineret af familien Angkatells sære opførsel, så han siger ja tak til at tilbringe weekenden på deres landsted. Opholdet bliver dog en del mere begivenhedsrigt, end den lille detektiv har forestillet sig. En af gæsterne findes skudt, og der er ikke mangel på mistænkte, for alle i huset havde et horn i siden på afdøde. Poirot: David Suchet. John Christow: Jonathan Cake. Gudgeon: Edward Fox. Lady Angkatell: Sarah Miles. Instruktion: Simon Langton. (t). Genre : Serier. Year : 1994
DR1|1463928300|Kriminalkommissær Barnaby (11)|||0|0||Engelsk krimiserie."En fremmeds død". Barnaby holder ferie, og i hans fravær arresterer hans kollega Pringle en ung krybskytte for mordet på en vagabond, der er fundet død i skoven efter en rævejagt. Barnaby har dog ikke megen tiltro til sin kollegas dømmekraft, og da det lille landsbysamfund rammes af endnu et mistænkeligt dødsfald, beslutter han sig for at genåbne sagen. (t). Episode : 11. Genre : Serier. Year : 1999
DR1|1463934600|TV AVISEN med Sporten|||0|0||TV AVISEN med Sporten
DR1|1463936700|Dyrebørnenes første tid (2:5)||2012|0|0||Naturserie fra BBC fra 2012.Maj er den sværeste måned at være løve i Masai Mara i Kenya. Der er langt tid til, at gnuerne vandrer forbi, og føden er sparsom. Den fem måneder gamle løveunge, Moja, kæmper sammen med sin mor for at overleve. De er alene og tilhører ikke nogen flok, og det gør dem meget sårbare. Løver i en stor flok kan samarbejde om at nedlægge større byttedyrsom bøfler, der kan give mad til mange i flere dage. Det kan Moja og hans mor ikke, men da regnen kommer, og græsset begynder at gro, bringer det også håb om overlevelse for den lille tapre familie. (t). Episode : 2:5. Genre : Dokumentar. Year : 2012
DR1|1463940000|Natportieren - The Night Manager (6:6)||2016|0|0||Engelsk thrillerserie fra 2016 efter en roman af John Le Carré. Roper tager til Cairo med sit hold for at lukke våbenaftalen. I Cairo møder Pine sin gamle fjende. Pine beslutter at satse alt for at gennemføre sin dobbelte hævnaktion. London lukker ned for støtten til Steadman og Burrs antikorruptionsprogram og mens Roper lægger sidste hånd på aftalen, slås Pine og Burr for at redde operationen med livet som indsats. Serien er uegnet for børn. Medvirkende: Hugh Laurie, Tom Hiddleston, Olivia Colman m.fl. Manuskript: David Farr. Instruktion: Susanne Bier. Produktion: The Ink Factory for BBC. (t). Episode : 6:6. Genre : Serier. Year : 2016
DR1|1463943600|TV AVISEN|||0|0||TV AVISEN
DR1|1463946000|Fodboldmagasinet||2016|0|0||Få det fulde overblik over Superligaen, når DR1 hver søndag blænder op for Fodboldmagasinet. Vi viser højdepunkter fra alle weekendens kampe og har gæster med i studiet, når der skal sættes ord på den seneste udvikling i den bedste danske fodboldrække. Derudover er der sidste nyt fra de store udenlandske fodboldligaer og de mest væsentlige nyheder fra den øvrige sportsverden. Vært: Peter Møller. (t). Genre : Sport. Year : 2016
DR1|1463947800|Kommissær George Gently (20)||2015|0|0||Engelsk krimiserie fra 2015.Nordøstengland, 1969. En prostitueret anmelder en voldtægt. Efterfølgende opdager kommissær Gently, at politiet har undladt at efterforske en lang række voldtægtssager. Den erfarne politimand er forfærdet og vil vide hvorfor. Sagen bliver ekstra presserende, da en kvinde findes voldtaget og myrdet. Nu går jagten på morderen ind. George Gently: Martin Shaw. John Bacchus: Lee Ingleby. Rachel Coles: Lisa McGrillis. Instruktion: Roger Goldby. (t). Episode : 20. Genre : Serier. Year : 2015
DR1|1463953200|30 grader i februar (5:10)||2012|0|0||<h2 class='program-small-desc'>Svensk dramaserie fra 2012Svensk dramaserie fra 2012.En række svenskere er taget til Thailand i jagten på et bedre liv. Krigen mellem de to Happiness Bungalows trappes op. Joy ved ikke, at Pong bor blot nogle få meter fra hende. Majlis har dræbt sin mand ved et uheld, og nu må hun finde ud af, hvad hun skal stille op med hans lig. Og Glenn møder Dits forældre. (t). Episode : 5:10. Genre : Film. Year : 1911
DR1|1463956500|Taggart: Mellem liv og død||2005|0|0||Skotsk krimiserie fra 2005.En fredelig fisketur udvikler sig dramatisk, da Matt Burke skydes ned af en ukendt gerningsmand. Samme dag bliver en politimand fra bedrageriafdelingen likvideret. I begges hjem finder efterforskningsholdet et stort pengebeløb i kontanter, og mens Burke kæmper for sit liv på hospitalet, må hans kolleger spørge sig selv, om deres chef har modtaget bestikkelse
DR1|1463960700|Amerikansk komediedrama fra 1987||1987|0|0||<h2 class='program-small-desc'>Amerikansk komediedrama fra 1987Amerikansk komediedrama fra 1987.Politimanden Burt Simpson erfarer, at han kun har kort tid tilbage at leve i. Burt beslutter sig for at blive dræbt på jobbet, så hans familie kan få udbetalt hans livsforsikring. Pludselig har stationen fået sig en ny superstrømer, der frygtløst kaster sig ud i de mest vanvittige situationer. Burt Simpson: Dabney Coleman. Ernie Dills: Matt Frewer. Carolyn: Teri Garr. Instruktion: Gregg Champion. (t). Genre : Film. Year : 1987
DR1|1463966100|Under Hammeren||2014|0|0||I Under Hammeren er alt på spil, når der rundt om i Danmark afholdes auktioner over alt fra blomster og kvæg til fine antikviteter og konkursboer. Hvem får solgt til prisen, og hvor langt er køberne egentlig villige til at gå. Følg med når auktionarius Kim Davidsen fra Sjællands Bilauktion sælger motorcykler for Politiet. Hos Thomas Rasmussen fra Blomsterauktionen Gasa skal en verdensnyhed under hammeren. Liselotte Møller fra Lauritz.com er på vurderingsbesøg hos Smartrooms, hvor der dukker flere usædvanlige møbler op. Sendt første gang 12.03.15 (t). Genre : Fritid & Livsstil. Year : 2014
DR1|1463967600|Kender Du Typen? (8:8)|||0|0||"Kender Du Typen?" er taget ud i sommerlandet, hvor en kendt dansker har indrettet sig i et sommerhus med værelse til svigermor og atelier til konen. Hvem er det, som er så vild med kvinderne i sit liv? Det skal livsstilseksperterne Anne Glad og Flemming Møldrup finde ud af i aftenens udsendelse. Vært: Mads Steffensen (t). Episode : 8:8. Genre : Fritid & Livsstil. Year : 2015
DR1|1463970300|Hammerslag (3)|||0|0||I aften er Hammerslag i Danmarks sydøstlige hjørne. Første stop er lidt udenfor Sakskøbing på Lolland. Hvad mon et sommerhus, en såkaldt flexbolig, koster på disse kanter? Aftenens anden bolig ligger i Hasselø på Falster, og er en kæmpevilla på mere end 300 m2. Det tog lang tid at sælge den, men hvad blev prisen? Vi slutter i Guldborg med en villa lige ud til vandet. Vil du gætte med på prisen? Se Hammerslag. Sendt første gang 16.09.14 (t). Episode : 3. Genre : Fritid & Livsstil. Year : 2014
DR1|1463977500|Overklassen på udebane (1:3)||2015|0|0||I Overklassen på udebane forlader modekongen Erik Brandt og dronningens tidligere ceremonimester, Christian Eugen-Olsen deres overklasseliv og bevæger sig ind i en ukendt verden, for at få sat ansigt på nogle af de mennesker, som de ellers kun hører om i statistikker og nyhedsindslag. I dag skal Erik og Christian besøge Annette Hansen fra Køge, der er enlig mor til tre og kassedame. Erik og Christian skal prøve at leve en dag i hendes liv, og mærke på egen krop, hvordan livet er udenfor deres privilegerede verden. 42-årige Annette er stolt af at være kassedame og blev i 2015 nomineret til at være årets sødeste kassedame. To grupper i samfundet, som sjældent møder hinanden, men kunne vi lære noget hvis vi gjorde. En morsom, rørende og nyskabende dokumentarserie på DR1 om ulighed. (t). Episode : 1:3. Genre : Dokumentar. Year : 2015
DR1|1463979300|De store katte (45)||1996|0|0||Naturserie fra BBC.Mød nogle af Kenyas mest karismatiske store katte i nationalparken Masai Mara. Her kæmper løver, geparder, og leoparder for at overleve i den storslåede, men ikke altid lige gæstfrie natur. (t). Episode : 45. Genre : Natur & Miljø. Year : 1996
DR1|1463981100|Verdens vildeste øer - Hebriderne (5:5)||2012|0|0||Hollandsk naturserie fra 2012.Verdens øer kan være hjemsted for nogle af de mest dramatiske landskaber og det mest fantastiske dyreliv. Mange tusinde års isolation har virket som brændstof på den naturlige udvælgelse, det vil sige tilpasningen til de særlige naturforhold, og har ikke alene fået de mest besynderlige væsner til at trives og overleve, men har også ført til en udvikling af nye arter specialiseret i at overleve de særlige naturforhold netop der. (t). Episode : 5:5. Genre : Natur & Miljø. Year : 2012
DR1|1463984100|De flyvende læger (184:224)|||0|0||Australsk dramaserie.I den lille australske flække Cooper's Crossing holder den flyvende lægetjeneste til. I den tyndt befolkede landsdel er der langt til lægen, så i stedet må læger og sygeplejersker flyve ud til områdets afsidesliggende gårde, kvægstationer og minelandsbyer for at yde lægehjælp - ofte under vanskelige og farlige forhold. (t). Episode : 184:224. Genre : Serier. Year : 1986
DR1|1463986800|De flyvende læger (185:224)|||0|0||Australsk dramaserie.I den lille australske flække Cooper's Crossing holder den flyvende lægetjeneste til. I den tyndt befolkede landsdel er der langt til lægen, så i stedet må læger og sygeplejersker flyve ud til områdets afsidesliggende gårde, kvægstationer og minelandsbyer for at yde lægehjælp - ofte under vanskelige og farlige forhold. (t). Episode : 185:224. Genre : Serier. Year : 1986
DR1|1463989500|Kystvagten (57:68)|||0|0||Australsk dramaserie.Narkosmugling, ulovligt fiskeri, menneskesmugling, ueksploderede miner og sågar terrorisme. Det er blot nogle af de problemer, der møder kaptajnløjtnant Mike Flynn og resten af besætningen på patruljebåden HMAS Hammersley, når de dagligt overvåger farvandet omkring Australiens kyster. Også blandt besætningen går bølgerne af og til højt. For det kan være sin sag at leve sammen i månedsvis på meget lidt plads. (t). Episode : 57:68. Genre : Serier. Year : 2007
DR1|1463991900|OBS|||0|0||Oplysning til borgerne om samfundet. (t). Genre : Forbruger. Year : 2016
DR1|1463992200|Antikkrejlerne (16)||2010|0|0||Britisk dokumentarserie fra 2010.Hver uge rejser to antikvitetseksperter med 200 pund på lommen til en egn af Storbritannien for i små antikvitetsbutikker at gå på jagt efter netop det fund, der kan indbringe køberen den største fortjenenste på den nærmeste auktion. (t). Episode : 16. Genre : Serier. Year : 2010
DR1|1463994000|Antikkrejlerne med kendisser (86)||2011|0|0||Britisk dokumentarserie fra 2011.Nogle af Storbritanniens kendteste antikvitetseksperter slår sig sammen med en række kendte i jagten på antikviteter og loppemarkedsfund. Hvilket hold kan skabe den største fortjeneste? (t). Episode : 86. Genre : Serier. Year : 2015
DR1|1463997600|Under Hammeren||2015|0|0||I Under Hammeren er alt på spil, når der rundt om i Danmark afholdes auktioner over alt fra blomster og kvæg til fine antikviteter og konkursboer. Hvem får solgt til prisen, og hvor langt er køberne egentlig villige til at gå. I dagens afsnit afholder Auktionshuset Hørsholm frimærkeauktion for første gang nogensinde. Hos Svendborg Auktion er der eftersyn, og så siges der også farvel til chefen gennem mange år, Jan Helmer. Og hos York Auktion har Ole Mortensen store forventninger til prisen på en gummibåd. (t). Genre : Fritid & Livsstil. Year : 2015
DR1|1463999400|Kender Du Typen? (1:10)|||0|0||Aftenens kendte hovedperson har skiftet storbylivet og caffe latterne ud med en tilværelse på landet og hjemmebrygget kaffe - og det har ikke været uden kultursammenstød. Det og meget mere lærer livsstilseksperterne Anne Glad og Flemming Møldrup om den hemmelige hovedperson, inden de til sidst skal regne ud, hvilken kendt dansker de er på besøg hos. Vært: Mads Steffensen (t). Episode : 1:10. Genre : Dokumentar. Year : 2016
DR1|1464001800|Hammerslag i Berlin|||0|0||Hammerslag er taget til Europas centrum, Berlin.Byen der har været bombet tilbage til stenalderen og derefter brutalt delt op af en mur i 30 år, har rejst sig igen. Danskerne køber lejligheder i Berlin for at leve livet på mærkelige cafeer og føle historiens vingesus i verdensbyen. Og så er det billigt at købe sig en bolig i storbyen - indtil videre. Hammerslag er udvidet til en time, så udover at gætte priser på boliger får du også en guide til alt det der gør Berlin til noget helt særligt. Østholdet. Ejendomsmægler Anders Gerner Frost og. ejendomsmægler Kristina Beck Poulsen. Vestholdet. Ejendomsmægler Claus Dreyer og. ejendomsmægler Inge Ørtoft. www.dr.dk/hammerslag. Sendt første gang 21.12.07 (t). Genre : Fritid & Livsstil. Year : 2007
DR1|1464005400|Johan Falk: GSI - Gruppen for særlige indsatser||2009|0|0||Svensk thriller fra 2009.I fem år har Johan Falk arbejdet for Europol i Haag. Nu vender han hjem til Göteborg, hvor han har fået job i politienheden GSI, der bekæmper grov organiseret kriminalitet. Her kastes Johan direkte ind i en risikofyldt operation, der går ud på at identificere og pågribe en brutal bande, der står bag en række voldsomme røverier mod pengetransporter. Johan Falk: Jakob Eklund. Frank Wagner: Joel Kinnaman. Patrik Agrell: Mikael Tornving. Instruktion: Anders Nilsson. (t). Genre : Serier. Year : 2010
DR1|1464012300|Taggart: Blodpenge||2002|0|0||Skotsk krimi fra 2002.Burke, Ross og Fraser har ringside-pladser, da bokseren Andy Corbett overraskende besejrer favoritten Jimmy Sullivan. Noget tyder på, at det er aftalt spil, og da kampens promoter findes dræbt, vender Burke søgelyset mod en gammel bekendt. For hvad har bragt gangsteren Sammy Cassidy hjem til Glasgow efter 20 år i USA. Jackie Reid: Blythe Duff. Robbie Ross: John Michie. Matt Burke: Alex Norton. Instruktion: Brian Kelly. (t). Genre : Serier. Year : 1996
DR1|1464015300|Jordemoderen IV (4:10)||2014|0|0||Engelsk dramaserie fra 2014.Londons East End, 1959. Med tilknytning til et nonnekloster hjælper en gruppe jordemødre, sygeplejersker og nonner den fattige bydels gravide kvinder. (t). Episode : 4:10. Genre : Serier. Year : 2014
DR1|1464018600|TV AVISEN|||0|0||TV AVISEN
DR1|1464019200|Under Hammeren||2015|0|0||I Under Hammeren er alt på spil, når der rundt om i Danmark afholdes auktioner over alt fra blomster og kvæg til fine antikviteter og konkursboer. Hvem får solgt til prisen, og hvor langt er køberne egentlig villige til at gå. I dagens afsnit afholder York Auktion eftersyn, og det tiltrækker flere mennesker end ventet, så Ole må holde nerverne i ro med en gammel vane. Hos Bruun Rasmussen sælges en yderst sjælden Poul Kjærholm-daybed, som Liselotte Toxværd Møller har store forventninger til. Og hos Sjællands Bilauktion har Kim Davidsen tre toiletvogne under hammeren, som viser sig at være ret eftertragtet. (t). Genre : Fritid & Livsstil. Year : 2015
DR1|1464021000|TV AVISEN med Sporten|||0|0||TV AVISEN med Sporten
DR1|1464022500|Vores vejr|||0|0||Vores vejr
DR1|1464023100|Aftenshowet||2016|0|0||DR1s journalistiske talkshow direkte fra Rådhuspladsen i København. (t). Genre : Underholdning. Year : 2016
DR1|1464026100|TV AVISEN|||0|0||TV AVISEN
DR1|1464026400|Bag Verden - med Tobias (3:6)|||0|0||Belgien.Tobias Hamann-Pedersen rejser til Belgien, som er en sværvægter inden for lækre delikatesser. Her bliver han blandt andet udfordret til at sniffe den verdensberømte belgiske chokolade og cykle hen over Belgiens berygtede brosten. Men landets høje standard inden for søde sager giver Tobias sved på panden, når han skal samle alle oplevelserne i én kage til sine belgiske værter. (t). Episode : 3:6. Genre : Ukategoriseret. Year : 2015
DR1|1464029100|En syg forskel (1:4)||2016|0|0||Jan har risiko for at dø tidligt. Han er arbejdsløs og bor i et socialt boligbyggeri i Aalborg. 7 kilometer derfra i et velhavende villakvarter lever de jævnaldrende mænd i snit 16 år længere end Jan. Hvorfor bliver nogle mere syge end andre? Er der forskel på den behandling rige og fattige får på hospitalet og hos lægen? I en ny serie undersøger DR Dokumentar uligheden i det danske sundhedssystem. Tilrettelæggelse: Lisbeth Dilling og Nikolaj Venge (t). Episode : 1:4. Genre : Dokumentar. Year : 2016
DR1|1464031800|TV AVISEN|||0|0||TV AVISEN
DR1|1464033300|Horisont|||0|0||Horisont
DR1|1464034800|Sporten|||0|0||Sporten
DR1|1464035400|Kriminalinspektør Banks: Begravet||2015|0|0||Engelsk krimi fra 2015.Liget af en fremtrædende kvindelig advokat skylles op på bredden af en underjordisk flod. Alan Banks får mistanke om, at morderen skal findes blandt medlemmerne af kvindens egen familie. Snart bliver der begået endnu et mord, og Banks må optrevle et net af hemmeligheder og løgne for at finde frem til gerningsmanden. Alan Banks: Stephen Tompkinson. Annie Cabbot: Andrea Lowe. Helen Morton: Caroline Catz. (t). Genre : Serier. Year : 2014
DR1|1464040800|Til undsætning (43:48)||2010|0|0||Australsk dramaserie fra 2010.De sætter livet på spil for at redde andre. De ansatte i den australske redningstjeneste Rescue Special Ops er nemlig eksperter i redningsmissioner af enhver art - til lands, til vands og i luften(n)
DR1|1464043500|To sønner (1:22)|||0|0||Amerikansk dramaserie.Mordet på Tom efterlader hans barnløse bror Rudy med to viljestærke sønner. Toms søn Wesley vokser op som en uregerlig kostskoleelev, mens Julies søn Billy udfolder sig som helikopterskytte i Vietnam(n)
DR1|1464046200|Kystvagten (1:68)|||0|0||Australsk dramaserie.Narkosmugling, ulovligt fiskeri, menneskesmugling, ueksploderede miner og sågar terrorisme. Det er blot nogle af de problemer, der møder kaptajnløjtnant Mike Flynn og resten af besætningen på patruljebåden HMAS Hammersley, når de dagligt overvåger farvandet omkring Australiens kyster. Også blandt besætningen går bølgerne af og til højt. For det kan være sin sag at leve sammen i månedsvis på meget lidt plads. Episode : 1:68. Genre : Serier. Year : 2007(n)
DR1|1464048900|Under Hammeren||2015|0|0||I Under Hammeren er alt på spil, når der rundt om i Danmark afholdes auktioner over alt fra blomster og kvæg til fine antikviteter og konkursboer. Hvem får solgt til prisen, og hvor langt er køberne egentlig villige til at gå. I dagens afsnit afholder Auktionshuset Hørsholm frimærkeauktion for første gang nogensinde. Hos Svendborg Auktion er der eftersyn, og så siges der også farvel til chefen gennem mange år, Jan Helmer. Og hos York Auktion har Ole Mortensen store forventninger til prisen på en gummibåd. Genre : Fritid & Livsstil. Year : 2015(n)
DR1|1464050700|Kender Du Typen? (1:10)|||0|0||Aftenens kendte hovedperson har skiftet storbylivet og caffe latterne ud med en tilværelse på landet og hjemmebrygget kaffe - og det har ikke været uden kultursammenstød. Det og meget mere lærer livsstilseksperterne Anne Glad og Flemming Møldrup om den hemmelige hovedperson, inden de til sidst skal regne ud, hvilken kendt dansker de er på besøg hos. Vært: Mads Steffensen. Episode : 1:10. Genre : Dokumentar. Year : 2016(n)
DR1|1464053400|Hammerslag i Berlin|||0|0||Hammerslag er taget til Europas centrum, Berlin.Byen der har været bombet tilbage til stenalderen og derefter brutalt delt op af en mur i 30 år, har rejst sig igen. Danskerne køber lejligheder i Berlin for at leve livet på mærkelige cafeer og føle historiens vingesus i verdensbyen. Og så er det billigt at købe sig en bolig i storbyen - indtil videre. Hammerslag er udvidet til en time, så udover at gætte priser på boliger får du også en guide til alt det der gør Berlin til noget helt særligt. Østholdet. Ejendomsmægler Anders Gerner Frost og. ejendomsmægler Kristina Beck Poulsen. Vestholdet. Ejendomsmægler Claus Dreyer og. ejendomsmægler Inge Ørtoft. www.dr.dk/hammerslag. Sendt første gang 21.12.07. Genre : Fritid & Livsstil. Year : 2007(n)
DR1|1464056700|70'erne tur retur: 1979|||0|0||Velkommen til 1970'ernes allersidste kapitel. I 1979 er der både håb og frygt for hvad fremtiden byder på. Genre : Ukategoriseret. Year : 2013(n)
DR1|1464063900|Overklassen på udebane (2:3)||2015|0|0||Modekongen Erik Brandt og den tidligere ceremonimester Christian Eugen-Olsen er virkelig på udebane, når de besøger en ung arbejdsløs kvinde, som bor i en lejlighed på et værelse i Albertslund. Langt væk fra Strandvejen og Eriks 400 kvadratmeter store herskabslejlighed i København K. Heidi på 28 år er en af de mange unge i Danmark, som er ramt af arbejdsløshed. Hun kæmper hver dag for at få et job. I dag skal Heidi og de to fine herre i virksomhedspraktik som stuepiger på et fint hotel i København. Heidi håber på at kunne imponere oldfruen, så hun vil kunne få et job på hotellet, når de skal ansætte nye stuepiger. Erik og Christian kæmper for at følge med Heidi, men det er tydeligt, at de ikke selv er vant til at stå for rengøringen derhjemme. Som Erik siger: 'Jeg har ikke redt min egen seng i 50 år.'.OVERKLASSEN PÅ UDEBANE er en sjov og tankevækkende serie om ulighed i Danmark. Episode : 2:3. Genre : Dokumentar. Year : 2015(n)
DR1|1464065700|De store katte (46)||1996|0|0||Naturserie fra BBC.Mød nogle af Kenyas mest karismatiske store katte i nationalparken Masai Mara. Her kæmper løver, geparder, og leoparder for at overleve i den storslåede, men ikke altid lige gæstfrie natur. Episode : 46. Genre : Natur & Miljø. Year : 1996(n)
DR1|1464067500|Vilde fødsler - Elefanter||2015|0|0||Britisk naturserie fra 2015.Dyrlægen Mark Evans og anatomen Joy Reidenberg udforsker de vidunderlige og ind imellem temmelig mærkværdige måder, som dyr føder deres unger på. Først besøger de Afrika for at undersøge de specielle vanskeligheder, som jordens største landdyr, elefanten, står over for, når den skal forplante sig og føde sunde unger. Genre : Dokumentar. Year : 2015(n)
DR1|1464070500|De flyvende læger (186:224)|||0|0||Australsk dramaserie.I den lille australske flække Cooper's Crossing holder den flyvende lægetjeneste til. I den tyndt befolkede landsdel er der langt til lægen, så i stedet må læger og sygeplejersker flyve ud til områdets afsidesliggende gårde, kvægstationer og minelandsbyer for at yde lægehjælp - ofte under vanskelige og farlige forhold. Episode : 186:224. Genre : Serier. Year : 1986(n)
DR1|1464073200|De flyvende læger (187:224)|||0|0||Australsk dramaserie.I den lille australske flække Cooper's Crossing holder den flyvende lægetjeneste til. I den tyndt befolkede landsdel er der langt til lægen, så i stedet må læger og sygeplejersker flyve ud til områdets afsidesliggende gårde, kvægstationer og minelandsbyer for at yde lægehjælp - ofte under vanskelige og farlige forhold. Episode : 187:224. Genre : Serier. Year : 1986(n)
DR1|1464075900|Kystvagten (58:68)|||0|0||Australsk dramaserie.Narkosmugling, ulovligt fiskeri, menneskesmugling, ueksploderede miner og sågar terrorisme. Det er blot nogle af de problemer, der møder kaptajnløjtnant Mike Flynn og resten af besætningen på patruljebåden HMAS Hammersley, når de dagligt overvåger farvandet omkring Australiens kyster. Også blandt besætningen går bølgerne af og til højt. For det kan være sin sag at leve sammen i månedsvis på meget lidt plads. Episode : 58:68. Genre : Serier. Year : 2007(n)
DR1|1464078300|Antikkrejlerne (17)||2010|0|0||Britisk dokumentarserie fra 2010.Hver uge rejser to antikvitetseksperter med 200 pund på lommen til en egn af Storbritannien for i små antikvitetsbutikker at gå på jagt efter netop det fund, der kan indbringe køberen den største fortjenenste på den nærmeste auktion. Episode : 17. Genre : Serier. Year : 2010(n)
DR1|1464080100|Antikkrejlerne med kendisser (87)||2011|0|0||Britisk dokumentarserie fra 2011.Nogle af Storbritanniens kendteste antikvitetseksperter slår sig sammen med en række kendte i jagten på antikviteter og loppemarkedsfund. Hvilket hold kan skabe den største fortjeneste. Episode : 87. Genre : Serier. Year : 2015(n)
DR1|1464083700|Under Hammeren||2015|0|0||I Under Hammeren er alt på spil, når der rundt om i Danmark afholdes auktioner over alt fra blomster og kvæg til fine antikviteter og konkursboer. Hvem får solgt til prisen, og hvor langt er køberne egentlig villige til at gå. I dagens afsnit ankommer der ekstra mange dyr til Aars Landboauktion, så der er kamp om pladserne. Hos Sjællands Bilauktion skal Kim Davidsen sælge en bil, man ikke ser hver dag. Og i Svendborg er det Jan Helmers sidste dag som ejer af Svendborg Auktionerne. Genre : Fritid & Livsstil. Year : 2015(n)
DR1|1464085500|Kender Du Typen? (2:10)|||0|0||Hvilken kendt dansker taler til sin stuebirk, vasker sine gummisko med speciel shampoo og elsker hot sauce? Det skal livsstilseksperterne Anne Glad og Flemming Møldrup finde ud af, når de tager på opdagelse i en stor, nyrenoveret lejlighed på Nørrebro. Vært: Mads Steffensen. Episode : 2:10. Genre : Fritid & Livsstil. Year : 2016(n)
DR1|1464087900|Hammerslag Sommermix (4:4)||2012|0|0||Peter Ingemann har fundet de bedste, sjoveste, skæveste, dyreste, billigste og mest interessante boliger fra de sidste 8 år. Der bliver vist klip fra før, under og efter finanskrisen, og der bliver fortalt historier fra programmet - også når kameraerne er slukket. Sendt første gang 17.07.12. Episode : 4:4. Genre : Fritid & Livsstil. Year : 2012(n)
DR1|1464089700|Johan Falk: Våbenbrødre||2009|0|0||Svensk thriller fra 2009.Johan Falk har fået job i specialenheden GSI, der bekæmper grov organiseret kriminalitet. En rutineopgave afslører, at nogen i Göteborgs underverden er ved at samle våben nok til en mindre krig. Johan håber, at hans meddeler Frank Wagner kan skaffe oplysninger, der kan afsløre, hvad der foregår. Men for Frank bliver sagen et mareridt, da det går op for bandelederen Seth, at der er en stikker blandt hans folk. Johan Falk: Jakob Eklund. Frank Wagner: Joel Kinnaman. Asim Popov: Thomas W. Gabrielsson. Instruktion: Anders Nilsson. Genre : Serier. Year : 2010(n)
DR1|1464095400|Bergerac: Kærestesorger||1991|0|0||Engelsk krimi fra 1991.Danielle slår op med Jim Bergerac, der forsøger at drukne sine sorger på bunden af en flaske. Charlie er. bekymret for sin ven, og hans løsning er at holde Bergerac beskæftiget. Han overtaler ham til at tage med til. byen Bath for at passe på et værdifuldt maleri. Her lader den kærlighedssyge eksstrømer sig forblinde af en smuk kvinde, der absolut ikke har reelle hensigter. Genre : Serier. Year : 2003(n)
DR1|1464101700|Jordemoderen IV (5:10)||2015|0|0||Engelsk dramaserie fra 2015.Londons East End, omkring 1960. Med tilknytning til et nonnekloster hjælper en gruppe jordemødre, sygeplejersker og nonner den fattige bydels gravide kvinder. Episode : 5:10. Genre : Serier. Year : 2014(n)
DR1|1464105000|TV AVISEN|||0|0||TV AVISEN(n)
DR1|1464105600|Under Hammeren||2015|0|0||I Under Hammeren er alt på spil, når der rundt om i Danmark afholdes auktioner over alt fra blomster og kvæg til fine antikviteter og konkursboer. Hvem får solgt til prisen, og hvor langt er køberne egentlig villige til at gå. I dagens afsnit håber Heidi og Rikke fra Horsens Auktioner, at særligt et helt nummer vil lokke kunderne til eftersyn. Hos Dansk Maskinbørs kæmper Johannes med at presse priserne i vejret. Og hos Svendborg Auktionerne tester auktionarius Martin Nielsen et nyt system i håb om at lokke kineserne til at byde på et par fine vaser. Genre : Fritid & Livsstil. Year : 2015(n)
DR1|1464107400|TV AVISEN med Sporten|||0|0||TV AVISEN med Sporten(n)
DR1|1464108900|Vores vejr|||0|0||Vores vejr(n)
DR1|1464109500|Aftenshowet||2016|0|0||DR1s journalistiske talkshow direkte fra Rådhuspladsen i København. Genre : Underholdning. Year : 2016(n)
DR1|1464112500|TV AVISEN|||0|0||TV AVISEN(n)
DR1|1464112800|Kære nabo - gør bras til bolig - Frederiksberg|||0|0||Da Mai og Lars Serup mødte hinanden, boede Lars alene i en rummelig lejlighed på Frederiksberg - kun i selskab med sin 2-årige datter, Olivia, der boede der sammen med ham på halv tid. Og da Mai kort efter flyttede sine sparsomme Ikeamøbler ind i lejligheden, gjorde de ikke det store nummer ud af indretningen - det var de alt for forelskede til at tænke på. Seks år og to børn senere er Mai og Lars ved at drukne i bastante møbler, børnene har ikke plads til at lege på deres deleværelse - og familien lever af to gange SU og Lars' fritidsjob. Det halter med andre ord faktisk noget med både økonomi og overskud, og derfor har familien skrevet til designer, Natalia Sanchez, og skattejæger, Søren Falk, for at bede om hjælp. Og hjælp får de, når Kære Nabo-holdet og en flok gode naboer i andelsforeningen forbarmer sig over dem og tryller med gode genbrugsfund og masser af knofedt. Genre : Fritid & Livsstil. Year : 2016(n)
DR1|1464115500|Aldrig for sent (2:4)||2015|0|0||Peter og Stefanie. Hver femte dansker har på grund af en konflikt mistet kontakten til et eller flere familiemedlemmer. Stefanie er 18 år og har ikke set sin far siden hun blev tvangsfjernet da hun var ca. 2 år. Nu skal de med hjælp fra psykolog og familieterapeut Ulla Dyrløv møde hinanden. Et møde der vil åbne op for fortiden og et møde der vil ende i en forsoning eller et farvel. Stefanie er vokset op i gode plejefamilier, og ser stadig sin mor, men ingen af dem synes det er en god ide at hun møder Peter. Det er aldrig for sent at give hinanden en chance til og nu vil Stefanie endelig møde sin far, for at finde ud af om han er det monster hun igennem hele sit liv har fået fortalt han er. Episode : 2:4. Genre : Dokumentar. Year : 2015(n)
DR1|1464118200|TV AVISEN|||0|0||TV AVISEN(n)
DR1|1464119700|Sundhedsmagasinet: Overgangsalder|||0|0||Alle kvinder kommer i overgangsalderen. I langt de fleste tilfælde kan symptomerne behandles medicinsk. Men nogle fødevarer kan også have stor effekt. Værter: Lillian Gjerulf Kretz og Peter Qvortrup Geisling. Genre : Sundhed & Mad. Year : 2016(n)
DR1|1464121200|Sporten|||0|0||Sporten(n)
DR1|1464121800|Johan Falk: Leo Gaut||2009|0|0||Svensk thriller fra 2009.En nådesløs krig om Göteborgs restauranter er blusset op, og da en restaurationsejers bil bliver sprængt i luften uden for en skole, sætter Johan Falk og GSI alt ind på at stoppe krigen. Sagen bringer Johan Falk i forbindelse med en gammel kending, nemlig Leo Gaut. Eksforbryderen Gaut er nu lovlydig restaurantejer - og under hårdt pres fra gangstere, der ønsker at overtage hans forretning. Johan Falk: Jakob Eklund. Leo Gaut: Peter Andersson. Helén: Marie Richardson. Instruktion: Richard Holm. Genre : Serier. Year : 2010(n)
DRRAMA|1463868000|Godnat - Ramasjang|||0|0||Godnat - Ramasjang(n)
DRRAMA|1463889600|Gæt med Emil|||0|0||Op og ned på vippen
DRRAMA|1463890200|Gurli Gris|||0|0||Skygger. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463890500|Nysgerrige Nille|||0|0||Frihed
DRRAMA|1463891400|Kate og Mim-Mim|||0|0||Fuld frø frem
DRRAMA|1463892300|Thomas og hans venner|||0|0||Dukkefilm med dansk tale.Om det lille damptog Thomas og hans venner
DRRAMA|1463893200|Peter Kanin|||0|0||Historien om fru Snadreands æg
DRRAMA|1463894100|F for får|||0|0||F for får
DRRAMA|1463895000|Peter Plys: Forår i Hundredemeterskoven|||0|0||Tegnefilm med dansk tale
DRRAMA|1463898900|Op og hop (6)|||0|0||Nu skal du Op og hop. Kig med ind i Ramasjangs gymnastiksal og se hvordan du får gang i kroppen. Det gælder om at have det sjovt og få bevæget sig en helt masse, når Ramasjangs værter finder på gode øvelser. Uanset om du står i din stue eller på dit værelse kan du være med. For værterne i Ramasjang vil have alle i gang. Denne gang med Onkel Reje, der viser hvad dyrene i Zoo laver om natten. Episode : 6. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1463899500|Gurli Gris|||0|0||Bedste Kanins Dinosaurpark. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463899800|Gurli Gris|||0|0||Godnathistorie. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463900100|Gurli Gris|||0|0||Tabte nøgler. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463900400|Paw Patrol|||0|0||Vestens vilde vovser. Genre : For de mindste. Year : 2014
DRRAMA|1463901900|Chuggington|||0|0||Fut-tog trækning
DRRAMA|1463902500|Chuggington|||0|0||Hodges flyvetur
DRRAMA|1463903100|Paphoved (6:8)|||0|0||Potobferne. Papper er et paphoved og har ingen venner. Allerhelst vil han være venner med Lena, den cooleste pige i verden. Og så er den sure vicevært efter ham, indtil Papper fortæller ham at de farlige Potobfer kommer. Episode : 6:8. Genre : Børn & Ungdom. Year : 2011
DRRAMA|1463903400|Friends|||0|0||Stephanies fødselsdag. Genre : For større børn. Year : 2013
DRRAMA|1463904600|Eventyrdetektiven Sandra|||0|0||Kaptajn Sortskæg
DRRAMA|1463905500|Eventyrdetektiven Sandra|||0|0||Vejviserens tjerner
DRRAMA|1463906400|Dora udforskeren|||0|0||Dora udforskeren
DRRAMA|1463908200|Vilde venner II (8)|||0|0||Der er altid travlt i Vilde Venners klub hvor børn redder og passer på Danmarks vilde dyr. I dag er det Aske og Ellen, der har vagten i klubhuset. Der er efterårsrengøring på basen, så dyreburerne skal renses og sikres mod regnen. Og så skal Vilde Venner hjælpe en ged, der er kommet langt væk hjemmefra. Episode : 8. Genre : Børn & Ungdom. Year : 2013
DRRAMA|1463909400|Postmand Per|||0|0||En besværlig transportDukkefilm. Det er snevejr i Grønnedal, og da postbilen bryder sammen, må Per ud at låne et køretøj. Men det lader til at være en dårlig dag for biler og motorcykler. Genre : For de mindste. Year : 2005
DRRAMA|1463910300|Bamses Billedbog|||0|0||Hvem skal passe Lunas bål. Genre : For de mindste. Year : 1995
DRRAMA|1463911800|Ellevilde Ella|||0|0||Bamsen BammeBamsen Bamme
DRRAMA|1463912400|Dyrene fra Lilleskoven (8:13)|||0|0||Som far, sådan sønnen.Modig er taget ud for at klare sig selv. Imens planlægger Ræv et angreb på Skramme, men det bliver alting kun værre af
DRRAMA|1463913900|Køkkenhyggen Hella|||0|0||Klipse klapse fangeren.Fisker Holm kommer på besøg med en spand fyldt med vand og hemmeligheder. Genre : For de mindste. Year : 2012
DRRAMA|1463915400|Eventyrdetektiven Sandra|||0|0||Eventyrdetektiven Sandra
DRRAMA|1463916000|Nysgerrige Nille|||0|0||Helt absurd, Nille
DRRAMA|1463916600|Skæg med Ord|||0|0||Hr. Skæg tager på eventyr i en verden af ord. Han bliver inviteret på skovtur et hemmeligt sted, og han prøver igen at få Ordklaveret til at virke. I købmandsbutikken prøver Fejedrengen Jas at hjælpe Hr. Skæg med at købe ind, og så møder Hr. Skæg et kækt lille dyr, som kan larme og synge med konsonanter. Genre : For de mindste. Year : 2012
DRRAMA|1463918400|Brandmand Sam|||0|0||En dag ved kysten. Genre : For de mindste. Year : 2008
DRRAMA|1463919000|Thomas og hans venner|||0|0||Dukkefilm med dansk tale.Om det lille damptog Thomas og hans venner
DRRAMA|1463919600|Musen Tip|||0|0||På job med far
DRRAMA|1463920200|Ring til Ramasjang|||0|0||Bamsen Holger står i lidt af et dilemma: Han leger kyssefange med de andre bamser, men han vil kun kysses af Trille. Hvad gør han? Lille Skille har også et problem, for han har klædt sig ud som spøgelse og er blevet bange for sit eget spejlbillede
DRRAMA|1463920800|Det mindste kongerige i verden (5)|||0|0||Hulen. I Det mindste kongerige i verden, har troldmanden Pokus og Kongen travlt med at lære Prinsesse Krinoline alt, hun skal lære, for at blive en god dronning. Det kan godt være lidt kedeligt, men da Krinoline flytter ud i skoven, og møder en hulemand, sker der endelig noget spændende. Episode : 5. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1463922300|Dora udforskeren|||0|0||Dora udforskeren
DRRAMA|1463923800|Lille NØRD|||0|0||Struds.Nu skal Lille Nørd på tur! Rosa og Johan kører ud og besøger bondegårdsdyr på deres seje tandem, og cykelvognen er spækket med overraskelser. Så skal der leges. Værter: Rosa Nyholm og Johan Sarauw. Genre : For de mindste. Year : 2007
DRRAMA|1463925600|Gurli Gris|||0|0||Den hemmelige klub. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463925900|Gurli Gris|||0|0||Bedste Kanins bådplads. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463926200|Smølferne|||0|0||Smølferne
DRRAMA|1463927700|Doktor McStuffins||2013|0|0||Doktor McStuffins er altid klar til at hjælpe bamser, dukker og andet legetøj, der ikke har det godt. Hun har nemlig forvandlet sit legehus til en lægeklinik, hvor hun behandler alt fra dehydrerede brandbiler til deprimerede dukker. For når Doktor McStuffins tager sit magiske stetoskop på, bliver hendes legetøj levende. Genre : For de mindste. Year : 2013
DRRAMA|1463929200|Det kongelige spektakel|||0|0||Det Kongelige Spektakel er havnet i klitterne - tæt på vandet i det halve kongerige
DRRAMA|1463930100|Ramajetterne|||0|0||Flummer driller. Der er travlhed i lufthavnen, og når selveste Onkel Reje skal ud at rejse, skal han naturligvis have VIP-behandling. Alle får spændende opgaver undtagen Flummer, der udtænker en drilsk plan. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1463931600|Da Lotte blev usynlig|||0|0||Andet afsnit i serien om den snart syv-årige Lotte. Hun har fået en underlig 'knap' på maven. Når man trykker på den, forsvinder hun. Lottes storebror Øffe øjner chancen for at tjene penge på Lottes helt specielle evner. Genre : For de mindste. Year : 1988
DRRAMA|1463933100|Tree Fu Tom|||0|0||En rutsjetur i hulenEn rutsjetur i hulen. Genre : For de mindste. Year : 2014
DRRAMA|1463934600|Min oldefars historier - Fisketuren|||0|0||FisketurenTheodor er 5 år. Han er på besøg hos sin eventyrlige og (u)hyggelige Oldefar, som bor på en bjergtop langt oppe i Norge sammen med den lille kat Bombi Bitt
DRRAMA|1463935200|Ring til Ramasjang|||0|0||Bamsen Holger står i lidt af et dilemma: Han leger kyssefange med de andre bamser, men han vil kun kysses af Trille. Hvad gør han? Lille Skille har også et problem, for han har klædt sig ud som spøgelse og er blevet bange for sit eget spejlbillede
DRRAMA|1463935800|Molevitten|||0|0||Få et godt grin med Molevitten. Maskinen er endnu en gang landet i børnehaven, hvor friske unger sender sjove ting direkte til Hr. Skæg, Øvst, Silja og alle vennerne i Ramasjang. For hver ting de sender, får de en skør sketch retur
DRRAMA|1463936400|Eventyrdetektiven Sandra|||0|0||Kæmpe kærlighed
DRRAMA|1463937300|Yakari|||0|0||Indianerdrengen Yakari har en fantastisk evne: Han kan tale med dyr. Men med sådan en gave følger også et stort ansvar, for han vil hjælpe alle naturens skabninger, store som små - og det fører til mange farefulde oplevelser. Genre : Børn & Ungdom. Year : 2005
DRRAMA|1463938200|Abevej 64|||0|0||Amandas naboer
DRRAMA|1463938800|Kate og Mim-Mim|||0|0||Fuld frø frem
DRRAMA|1463939400|Godnathistorier|||0|0||Det er blevet aften i Ramasjang og tid til at sige tak for i dag. Men før vi slukker lyset og siger godnat, er der lige tid til en rigtig go' godnathistorie. Hr. Skæg læser op af Cirkus Saragossa. Genre : Børn & Ungdom. Year : 2013
DRRAMA|1463940000|Godnat - Ramasjang|||0|0||Godnat - Ramasjang
DRRAMA|1463976000|Gæt med Emil|||0|0||Natursamling
DRRAMA|1463976600|Gurli Gris|||0|0||International dag. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1463976900|Nysgerrige Nille|||0|0||Fordomme
DRRAMA|1463977800|Lille Nørd|||0|0||Kan det virkelig passe, at en græshoppe spiser vorter? Tag med Lille Nørd på græshoppejagt, og se hvordan Katrine bliver reddet af en østrigsk mesterdirigent. Leg med Lille Nørd på dr.dk/oline. Genre : For de mindste. Year : 2009
DRRAMA|1463979600|Kriblekrable Safari i haven|||0|0||De små dyr er lige omkring os. I dag tager børnene på kriblekrable safari i hus og have, hvor der er fyldt med spændende dyr
DRRAMA|1463980200|MikroMakkerne - Krible Krable|||0|0||MikroMakkerne har pakket deres trækvogn og er rullet ud i naturen for at gå på krible krable-jagt. I dag er det myren, som Selma og Milton skal blive klogere på. Dyk med dem ned i myretuen og find ud af, hvor sej den lille fætter egentlig er. Genre : Ukategoriseret. Year : 2016
DRRAMA|1463980800|Krible Krable ved vandet|||0|0||Krible Krable i vandet.Silja Okking tager til Bovbjerg Fyr og går på jagt efter Krible Krable-dyr i vandet. Imens er Sebastian Klein ved at gøre klar til fredagens store fest for alle de små, seje dyr
DRRAMA|1463982600|Vilde Venner - Krible Krable (1:5)|||0|0||Der er altid travlt i Vilde Venners klub, og i dag er det Aske og Ellen, der har vagten i klubhuset. Dagen står i de små krible-krable-dyrs tegn, så de tager en tur ud til Bjørli, der bor i skoven. Der går de på jagt efter smådyr i skovbunden, og når de kommer tilbage, har Bjørli en stor overraskelse til dem i køkkenet. For kan man egentlig spise små dyr man finder i skoven. Episode : 1:5. Genre : Ukategoriseret. Year : 2014
DRRAMA|1463983200|Ring til Ramasjang|||0|0||I dette afsnit ringer Hundsen, fordi han er ked af det. De andre bamser gider ikke at lege med ham, og han ved ikke, hvad han skal gøre. Elefanten Gumle ringer også, fordi der er en myg inde på værelset, og han er lidt nervøs for, hvad den kan finde på
DRRAMA|1463983800|Det kongelige spektakel|||0|0||Det Kongelige Spektakel er havnet i klitterne - tæt på vandet i det halve kongerige
DRRAMA|1463984700|Ramajetterne|||0|0||Flummer driller. Der er travlhed i lufthavnen, og når selveste Onkel Reje skal ud at rejse, skal han naturligvis have VIP-behandling. Alle får spændende opgaver undtagen Flummer, der udtænker en drilsk plan. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1463986200|Tree Fu Tom|||0|0||Træffel TomTræffel Tom. Genre : For de mindste. Year : 2012
DRRAMA|1463987400|Monster Buster|||0|0||Esther er rigtigt træt at sit dumme fantasi-monster, der har flagermusevinger og masser af øjne. Heldigvis kommer MonsterBuster Silja med klæd-ud-tøj og nogle seje flagermusevinger, og sammen buster de Esthers monster langt væk. For selvom monstre ikke findes i virkeligheden, kan man godt være bange for dem - og have brug for hjælp til at få dem væk. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1463988300|Peter Kanin|||0|0||Historien om den mystiske blommetyv
DRRAMA|1463989200|Ramasjang Mysteriet||2013|0|0||Hvor er Skoleinspektørens maltbolsjer? Der sker mystiske ting i Ramasjang. Byens syv skurke driller, og ting forsvinder. Heldigvis har Kristian en hemmelig detektivhule under byen, hvor han med hjælp fra superseje børn løser dagens mysterium. Genre : Børn & Ungdom. Year : 2013
DRRAMA|1463991000|Babar|||0|0||Operation Hemmelig Byttehandel. Genre : Børn & Ungdom. Year : 2010
DRRAMA|1463991900|Skæg med tal|||0|0||Et sjovt tælleprogram for de mindste med musik, dyr og masser af børn. Mød Hr. Skæg, som er vild med tal og med sit flotte, lange skæg. Mød også Regitze i butikken hvor man kun kan få én af hver vare. Og tag med Hr. Skæg, når han besøger børnenes små hemmelige restauranter, hvor der serveres frække deller, skøre isdesserter og meget, meget mere. Genre : For de mindste. Year : 2007
DRRAMA|1463993100|Gæt med Emil|||0|0||Mariehøns
DRRAMA|1463993700|Gæt med Emil|||0|0||Lille fugl spiser salatfrøene
DRRAMA|1463994600|Vilde venner II (9)|||0|0||Der er altid travlt i Vilde Venners klub hvor børn redder og passer på Danmarks vilde dyr. I dag er det Otto og Kaja der har vagten i klubhuset. Dyrlægen kommer på besøg for at undersøge og kastrere en hjemløs ged, og der skal bygges huler til små egernunger. Og så skal Vilde Venner redde en svane, der har forvildet sig ind i en boligblok. Episode : 9. Genre : Børn & Ungdom. Year : 2013
DRRAMA|1463995800|Postmand Per|||0|0||TordenvejretDukkefilm. Fru Madsen er bange for tordenvejr, og det er Poul også. Men da Bonny bliver væk, må nogen jo ud at finde den. Og Poul melder sig frivilligt. Genre : For de mindste. Year : 2005
DRRAMA|1463996700|Bamses Billedbog|||0|0||Bamse Dyregod og Knud Kylling. Genre : For de mindste. Year : 1995
DRRAMA|1463998200|Ellevilde Ella|||0|0||KagekonkurrencenKagekonkurrencen
DRRAMA|1463998800|Dyrene fra Lilleskoven (9:13)|||0|0||På et hængende hår.Stakkels Modig får brug for sine nye venner udenfor parken. Og inde i parken raser krigen mellem de gamle ræve, mens deres unger hellere vil slutte fred
DRRAMA|1464000300|Køkkenhyggen Hella|||0|0||Fuglene skal plukkes og steges.Det er jagt tid og 6 konger kommer til fest på klosteret. Genre : For de mindste. Year : 2012
DRRAMA|1464001800|Eventyrdetektiven Sandra|||0|0||Broder Trold
DRRAMA|1464002700|Nysgerrige Nille|||0|0||Du er for lille
DRRAMA|1464003000|Skæg med Ord|||0|0||Verdens allerførste ordHr. Skæg tager på eventyr i en verden af ord. Han bliver inviteret på skovtur et hemmeligt sted, og han prøver igen at få Ordklaveret til at virke. I købmandsbutikken prøver Fejedrengen Jas at hjælpe Hr. Skæg med at købe ind, og så synger Hr. Skæg om Ordmoderen, som opfandt verdens allerførste ord. Genre : For de mindste. Year : 2012
DRRAMA|1464004800|Brandmand Sam|||0|0||Brandmand Sam
DRRAMA|1464005400|Thomas og hans venner|||0|0||Dukkefilm med dansk tale.Om det lille damptog Thomas og hans venner
DRRAMA|1464006000|Musen Tip|||0|0||Hvor er Teddy
DRRAMA|1464006600|Ring til Ramasjang|||0|0||I dette afsnit ringer Trille, fordi hun leger far, mor og børn med de andre bamser - men hvad skal babyen hedde? Musikbamse ringer også, for han har en masse slik, som Fnuller kigger lige lovligt sultent på. Hvad skal han gøre
DRRAMA|1464007200|Det mindste kongerige i verden (6)|||0|0||Festmiddag. I Det mindste kongerige i verden, har troldmanden Pokus og Kongen travlt med at lære Prinsesse Krinoline alt, hun skal lære, for at blive en god dronning. Det kan godt være lidt kedeligt, men da Krinoline pludseligt får en baronesse til festmiddag, sker der endelig noget spændende. Episode : 6. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1464008700|Dora udforskeren|||0|0||Dora udforskeren
DRRAMA|1464010200|Lille Nørd|||0|0||Hvilket dyr skal Rosa og Johan møde i dag og hvad finder de mon på i deres hemmelige hule?. Tag med når "LilleNØRD" cykler ud på nye eventyr. Spil Lille Nørd på www.dr.dk/oline. Sendt første gang 5.10.08. Genre : For de mindste. Year : 2008
DRRAMA|1464011700|Gurli Gris|||0|0||Ryst, rasle og slå. Genre : Børn & Ungdom. Year : 2008
DRRAMA|1464012000|Gurli Gris|||0|0||Mester Far Gris. Genre : Ukategoriseret. Year : 2008
DRRAMA|1464012600|Smølferne|||0|0||Smølferne
DRRAMA|1464013800|Chuggington|||0|0||Wilson tager fat
DRRAMA|1464014400|Eventyrdetektiven Sandra|||0|0||Prinsesse af søen
DRRAMA|1464015600|Hej Ramasjang|||0|0||Vi roder og hamrer. Vi larmer og griner. Kom udenfor og ha' det sjovt med os i Hej Ramasjang. Hvem er sejest? Den tissende myre eller edderkoppen med sit spind? Det kribler og krabler ude ved laden i dag, hvor Silja og Rosa kæmper om at være det sejeste insekt. Genre : Børn & Ungdom. Year : 2015
DRRAMA|1464015660|Rosa fra Rouladegade||2011|0|0||Sophus' bilkage.Hvem skal man spørge, hvis man gerne vil have hjælp til at overraske nogen med en kage? Rosa fra Rouladegade selvfølgelig. Og det er lige netop hvad Sophus gør. Han vil nemlig gerne bage en kage til sin bedstefar, der har arbejdet som mekaniker og har sit helt eget bilværksted hjemme i garagen. Rosa og Sophus forklæder sig som gadefejere og sniger sig hjem til bedste, for at finde ud af hvad kagen skal ligne, hvilken farve den skal have og hvad den skal smage af. Genre : Børn & Ungdom. Year : 2011
DRRAMA|1464017700|MikroMakkerne - Krible Krable|||0|0||MikroMakkerne har pakket deres trækvogn og er rullet ud i naturen for at gå på krible krable-jagt. I dag smider de sig på maven og fanger krabber i nettet. Kig med, når Milton og Selma tester om krabben er så sej, som de tror, den er. Genre : Ukategoriseret. Year : 2016
DRRAMA|1464018300|Vilde venner krible krable|||0|0||Der er altid travlt i Vilde Venners klub, og i dag er det Aske og Ellen, der har vagten i klubhuset. Dagen står i de små krible-krable-dyrs tegn, så de tager en tur ud til Bjørli i skoven. De leder efter smådyr, for i dag vil de undersøge, om skovens myrer og bænkebiddere vil bo i deres hjemmelavede huse
DRRAMA|1464018600|Kriblekrable Safari hos myrerne|||0|0||Børnene er nysgerrige på at se hvordan myrer bor, så de bygger deres eget myrehotel
DRRAMA|1464019200|Ring til Ramasjang|||0|0||Møffe ringer fordi han bliver holdt udenfor af de andre bamser. Stritte ringer også til Ramasjang, for hendes hår klør så mærkeligt - hvad kan det mon skyldes
DRRAMA|1464020100|F for får|||0|0||Trafikprop
DRRAMA|1464020700|Nysgerrige Nille|||0|0||Helt absurd, Nille
DRRAMA|1464021300|Ramasjang Mysteriet|||0|0||Jacinta og Rasmus vandpistolerEr det Fru Pudderkvast, Danse Staffan eller en helt tredje der har været på spil? Der er i hvert fald ballade i Ramasjang! Jacinta og Rasmus har nemlig fået stjålet deres vandpistoler! Heldigvis får Kristian hjælp af minidetektiven Brage, men mon de kan finde den rigtige skurk? Se med i Ramasjang Mysteriet. Genre : Børn & Ungdom. Year : 2016
DRRAMA|1464022800|Peter Kanin|||0|0||Historien om Joakim Fiskers musikalske eventyrHistorien om Joakim Fiskers musikalske eventyr
DRRAMA|1464023700|Yakari|||0|0||Indianerdrengen Yakari har en fantastisk evne: Han kan tale med dyr. Men med sådan en gave følger også et stort ansvar, for han vil hjælpe alle naturens skabninger, store som små - og det fører til mange farefulde oplevelser. Genre : Børn & Ungdom. Year : 2005
DRRAMA|1464024600|Abevej 64|||0|0||Kamæleonen Kasper
DRRAMA|1464025200|Kate og Mim-Mim|||0|0||Ballonballade
DRRAMA|1464025800|Godnathistorier|||0|0||Det er blevet aften i Ramasjang og tid til at sige tak for i dag. Men før vi slukker lyset og siger godnat, er der lige tid til en rigtig go' godnathistorie. Hr. Skæg læser op af Cirkus Saragossa. Genre : Børn & Ungdom. Year : 2013
DRRAMA|1464026400|Godnat - Ramasjang|||0|0||Godnat - Ramasjang
DRRAMA|1464062400|Gæt med Emil|||0|0||Bløde ferskner (t)(n)
DRRAMA|1464063000|Gurli Gris|||0|0||Regnvejrsdag-legen (t). Genre : Børn & Ungdom. Year : 2008(n)
DRRAMA|1464063300|Nysgerrige Nille|||0|0||Biologiprøven (t)(n)
DRRAMA|1464064200|Lille Nørd|||0|0||Kan det virkelig passe, at myg godt kan lide sure tæer? Tag med Lille Nørd på mygge-eventyr, og se om det er Katrine eller Anders som kan få flest myggestik. Leg med Lille Nørd på dr.dk/oline (t). Genre : For de mindste. Year : 2009(n)
DRRAMA|1464066000|Kriblekrable Safari på stranden|||0|0||Børnene har sat en krabbefælde i havet. Dagen efter tømmer de den på stranden og ser, at det ikke kun er krabber, der er blevet lokket i fælden. (t)(n)
DRRAMA|1464066600|MikroMakkerne - Krible Krable|||0|0||MikroMakkerne har pakket deres trækvogn og er rullet ud i naturen for at gå på krible krable-jagt. I dag er det vårfluelarven, der skal fanges og undersøges. Se med om rygtet taler sandt og vårfluelarven kan bygge et hus af perler? (t). Genre : Ukategoriseret. Year : 2016(n)
DRRAMA|1464066900|Krible Krable i skoven|||0|0||Krible Krable i skoven.Silja Okking tager til Roskilde og går på jagt efter Krible Krable-dyr i skoven. Imens er Sebastian Klein ved at gøre klar til fredagens store fest for alle de små, seje dyr(n)
DRRAMA|1464068700|Vilde Venner - Krible Krable (2:5)|||0|0||Der er altid travlt i Vilde Venners klub, og i dag er det Aske og Ellen, der har vagten i klubhuset. Dagen står i de små krible-krable-dyrs tegn, så de tager en tur ud til Bjørli i skoven. De går på jagt efter forskellige snegle, og så laver de flotte slæder til Vilde Venners store sneglevæddeløb. (t). Episode : 2:5. Genre : Ukategoriseret. Year : 2014(n)
DRRAMA|1464069300|Ring til Ramasjang|||0|0||Dukke Nanna har brug for hjælp. Fnuller har spurgt hende, om de skal være kærester, men hvad laver kærester egentlig? Lille Isbjørn ringer også til Ramasjang, for der er en bi på værelset, og han ryster af skræk. (t)(n)
DRRAMA|1464069900|Lillefinger|||0|0||Den døde biMyren og Lillefinger finder en død bi ude i bakkerne og vil begrave den. Men bliver uenige om, hvordan man gør til en begravelse. (t). Genre : For de mindste. Year : 2009(n)
DRRAMA|1464070200|Rosa fra Rouladegade||2011|0|0||Sophus' bilkage.Hvem skal man spørge, hvis man gerne vil have hjælp til at overraske nogen med en kage? Rosa fra Rouladegade selvfølgelig. Og det er lige netop hvad Sophus gør. Han vil nemlig gerne bage en kage til sin bedstefar, der har arbejdet som mekaniker og har sit helt eget bilværksted hjemme i garagen. Rosa og Sophus forklæder sig som gadefejere og sniger sig hjem til bedste, for at finde ud af hvad kagen skal ligne, hvilken farve den skal have og hvad den skal smage af. (t). Genre : Børn & Ungdom. Year : 2011(n)
DRRAMA|1464072000|Tree Fu Tom|||0|0||Den fantastiske rejseDen fantastiske rejse. (t). Genre : For de mindste. Year : 2012(n)
DRRAMA|1464073200|Monster Buster|||0|0||Tvillingerne Alaska og Østen har problemer med hvert sit fantasi-monster. Østen har en dum zombie, og Alaska har en heks, der halter. Heldigvis ved MonsterBuster Mille lige, hvad der skal gøres - og sammen laver de tre en snedig fælde med mudder, sjove snorkelyde og et fangenet. For selvom monstre ikke findes i virkeligheden, kan man godt være bange for dem - og have brug for hjælp til at få dem væk. (t). Genre : Børn & Ungdom. Year : 2015(n)
DRRAMA|1464074100|Gurli Gris|||0|0||Ryst, rasle og slå (t). Genre : Børn & Ungdom. Year : 2008(n)
DRRAMA|1464074400|Peter Kanin|||0|0||Historien om den gnavne ugle. (t)(n)
DRRAMA|1464075300|Ramasjang Mysteriet||2013|0|0||Hvor er Kyllings mundharmonika? Der sker mystiske ting i Ramasjang. Byens syv skurke driller, og ting forsvinder. Heldigvis har Kristian en hemmelig detektivhule under byen, hvor han med hjælp fra superseje børn løser dagens mysterium. (t). Genre : Børn & Ungdom. Year : 2013(n)
DRRAMA|1464077100|Babar|||0|0||Fu finder (t). Genre : Børn & Ungdom. Year : 2010(n)
DRRAMA|1464077700|Babar|||0|0||Nålehovedet (t). Genre : Børn & Ungdom. Year : 2010(n)
DRRAMA|1464078600|Skæg med tal|||0|0||Et sjovt tælleprogram for de mindste med musik, dyr og masser af børn. Mød Hr. Skæg, som er vild med tal og med sit flotte, lange skæg. Mød også Regitze i butikken hvor man kun kan få én af hver vare. Og tag med Hr. Skæg, når han besøger børnenes små hemmelige restauranter, hvor der serveres frække deller, skøre isdesserter og meget, meget mere. (t). Genre : For de mindste. Year : 2007(n)
DRRAMA|1464079800|Gæt med Emil|||0|0||Op og ned på vippen (t)(n)
DRRAMA|1464081000|Vilde venner II (10)|||0|0||Der er altid travlt i Vilde Venners klub hvor børn redder og passer på Danmarks vilde dyr. I dag er det Otto og Kaja, der har vagten i klubhuset. Det nye ællingehus skal males, og der skal laves et rigtigt dejligt vinterbo til en skrubtudse. Og så skal Vilde Venner redde en fiskehejre, der er fanget i en fiskeline. (t). Episode : 10. Genre : Børn & Ungdom. Year : 2013(n)
DRRAMA|1464082200|Postmand Per|||0|0||Dr. Grøns fødselsdagsgaveDukkefilm. Per og Teddy vil gerne forære Dr. Grøn en bil, så hun lettere kan komme rundt til sine patienter, men hvor finder man lige en ledig bil? (t). Genre : For de mindste. Year : 2005(n)
DRRAMA|1464083100|Bamses Billedbog|||0|0||Ælling lærer at sige et ord. (t). Genre : For de mindste. Year : 1995(n)
DRRAMA|1464084600|Ellevilde Ella|||0|0||Orange dagOrange dag. (t)(n)
DRRAMA|1464085200|Dyrene fra Lilleskoven (10:13)|||0|0||Grævlings farvel.Væsel bliver anklaget og dømt for at stå i ledtog med Skramme. Og gamle Grævling tænker sig tilbage til sin lykkelige barndom i Lilleskoven, før han dør. I mellemtiden møder Modig en smuk hunræv i byen. (t)(n)
DRRAMA|1464086700|Køkkenhyggen Hella|||0|0||Næsten brækket ben og mexicansk mad.Storm og Emilie overrasker med indkøbsposer og aftensmad. (t). Genre : For de mindste. Year : 2012(n)
DRRAMA|1464088200|Eventyrdetektiven Sandra|||0|0||Scolymus (t)(n)
DRRAMA|1464088800|Nysgerrige Nille|||0|0||Frihed! (t)(n)
DRRAMA|1464089400|Skæg med Ord|||0|0||Hr. Skæg tager på eventyr i en verden af ord. Han bliver inviteret på skovtur et hemmeligt sted, og han prøver igen at få Ordklaveret til at virke. I købmandsbutikken prøver Fejedrengen Jas at hjælpe Hr. Skæg med at købe ind, og så synger Hr. Skæg om det ensomme bogstav K, som heldigvis møder O og R. (t). Genre : For de mindste. Year : 2012(n)
DRRAMA|1464091200|Brandmand Sam|||0|0||Brandmand Sam(n)
DRRAMA|1464091800|Thomas og hans venner|||0|0||Dukkefilm med dansk tale.Om det lille damptog Thomas og hans venner. (t)(n)
DRRAMA|1464092400|Musen Tip|||0|0||Jeg skal ikke til lægen (t)(n)
DRRAMA|1464093000|Ring til Ramasjang|||0|0||I dette afsnit ringer Fnuller, fordi han er i tvivl om, hvor meget slik, man egentlig kan spise uden at få ondt i maven. Snehvid ringer også. Han har brug for tips til at bygge en rigtig god hule. (t)(n)
DRRAMA|1464093600|Det mindste kongerige i verden (7)|||0|0||Portræt. I Det mindste kongerige i verden, har troldmanden Pokus og Kongen travlt med at lære Prinsesse Krinoline alt, hun skal lære, for at blive en god dronning. Det kan godt være lidt kedeligt, men da Krinoline skal have malet sit portræt af en kunstmaler, sker der endelig noget spændende. (t). Episode : 7. Genre : Børn & Ungdom. Year : 2015(n)
DRRAMA|1464095100|Dora udforskeren|||0|0||Dora udforskeren(n)
DRRAMA|1464096600|Lille Nørd|||0|0||Hvilket dyr skal Rosa og Johan møde i dag og hvad finder de mon på i deres hemmelige hule?. Tag med når "LilleNØRD" cykler ud på nye eventyr. Spil Lille Nørd på www.dr.dk/oline. Sendt første gang 21.10.08. (t). Genre : For de mindste. Year : 2008(n)
DRRAMA|1464098100|Gurli Gris|||0|0||Sludrechatol (t). Genre : Børn & Ungdom. Year : 2008(n)
DRRAMA|1464098400|Gurli Gris|||0|0||Hr. Rævs varevogn (t). Genre : Ukategoriseret. Year : 2008(n)
DRRAMA|1464099000|Smølferne|||0|0||Smølferne(n)
DRRAMA|1464100200|Chuggington|||0|0||Wilson og dinosaurussen (t)(n)
DRRAMA|1464100800|Eventyrdetektiven Sandra|||0|0||En uforglemmelig rejse (t)(n)
DRRAMA|1464102000|Hej Ramasjang|||0|0||Vi roder og hamrer. Vi larmer og griner. Kom udenfor og ha' det sjovt med os i Hej Ramasjang. Silja og Rosa kribler og krabler ude ved laden i dag. (t). Genre : Børn & Ungdom. Year : 2015(n)
DRRAMA|1464102060|Vilde venner II (8)|||0|0||Der er altid travlt i Vilde Venners klub hvor børn redder og passer på Danmarks vilde dyr. I dag er det Aske og Ellen, der har vagten i klubhuset. Der er efterårsrengøring på basen, så dyreburerne skal renses og sikres mod regnen. Og så skal Vilde Venner hjælpe en ged, der er kommet langt væk hjemmefra. (t). Episode : 8. Genre : Børn & Ungdom. Year : 2013(n)
DRRAMA|1464103500|Peddersen og Findus|||0|0||Peddersens telttur.Findus skal sove i telt - Alene! Det tør han alligevel ikke(n)
DRRAMA|1464104400|MikroMakkerne - Krible Krable|||0|0||MikroMakkerne har pakket deres trækvogn og er rullet ud i naturen for at gå på krible krable-jagt. I dag er det bænkebidderen, der bliver studeret nøje af Selma og Milton. Se med og bliv klogere på den lille grå fyr. (t). Genre : Ukategoriseret. Year : 2016(n)
DRRAMA|1464105000|Vilde venner krible krable|||0|0||Der er altid travlt i Vilde Venners klub, og i dag er det Asta og Sune, der har vagten i klubhuset. Dagen står i de små krible-krable-dyrs tegn, så de tager en tur ud til Bjørli i skoven. De tager på jagt efter smådyr i skoven, for Vilde Venner vil finde ud af, hvilket dyr, der er skovbundens hurtigste. (t)(n)
DRRAMA|1464105300|Kriblekrable Safari sommerfugle|||0|0||Der er både dag- og natsommerfugle, børnene sætter en lysfælde så de kan fange natsommerfugle, men de skal være hurtige, for fuglene vil gerne spise deres fangst. (t)(n)
DRRAMA|1464105900|Ring til Ramasjang|||0|0||I dette afsnit dratter Pelsi ned i håndvasken og bliver gennemblødt. Bamsen Pelle er ude på ballade - han har tænkt sig at lægge insekter i Fru Goks seng for at skræmme hende! (t)(n)
DRRAMA|1464106800|F for får|||0|0||Fårehyrden (t)(n)
DRRAMA|1464107400|Op og hop (10)|||0|0||Nu skal du Op og hop. Kig med ind i Ramasjangs gymnastiksal og se hvordan du får gang i kroppen. Det gælder om at have det sjovt og få bevæget sig en helt masse, når Ramasjangs værter finder på gode øvelser. Uanset om du står i din stue eller på dit værelse kan du være med. For værterne i Ramasjang vil have alle i gang. Denne gang med MonsterBuster der viser, hvordan de varmer op til at buste monstre. (t). Episode : 10. Genre : Børn & Ungdom. Year : 2015(n)
DRRAMA|1464108000|Dansebørnene i Cirkus Summarum 3:3||2015|0|0||Mød de seje dansebørn fra Cirkus Summarum. I dag er det den store premieredag. Alle er spændte! Nu skal dansebørnene og alle de andre i cirkus vise publikum det, de har øvet sig på. (t)(n)
DRRAMA|1464108900|F for får|||0|0||Den stinkende landmand (t)(n)
DRRAMA|1464109200|Peter Kanin|||0|0||Historien om det pibende legetøjHistorien om det pibende legetøj. (t)(n)
DRRAMA|1464110100|Yakari|||0|0||Indianerdrengen Yakari har en fantastisk evne: Han kan tale med dyr. Men med sådan en gave følger også et stort ansvar, for han vil hjælpe alle naturens skabninger, store som små - og det fører til mange farefulde oplevelser. (t). Genre : Børn & Ungdom. Year : 2005(n)
DRRAMA|1464110700|Abevej 64|||0|0||Simon Stork (t)(n)
DRRAMA|1464111600|Kate og Mim-Mim|||0|0||Glitrende Glimte. (t)(n)
DRRAMA|1464112200|Godnathistorier|||0|0||Det er blevet aften i Ramasjang og tid til at sige tak for i dag. Men før vi slukker lyset og siger godnat, er der lige tid til en rigtig go' godnathistorie. Hr. Skæg læser op af Cirkus Saragossa. (t). Genre : Børn & Ungdom. Year : 2013(n)
DRRAMA|1464112800|Godnat - Ramasjang|||0|0||Godnat - Ramasjang(n)
BBC Red Button 1|1463893200|FA Cup Football|FA Cup Goals: 2015/16 Final||0|0|Football - Club|Action from the final of the famous cup competition, as Crystal Palace faced Manchester United.
BBC Red Button 1|1463893200|FA Cup Football|FA Cup Goals: 2015/16 Final||0|0|Football - Club|Action from the final of the famous cup competition, as Crystal Palace faced Manchester United.
BBC Red Button 1|1463945100|EastEnders: Bobby: The Story So Far|||0|0|Soap,Melodrama|
BBC Red Button 1|1463979600|Mastertapes with Rufus Wainwright|Mastertapes: Paul McCartney||0|0|General Music,Ballet,Dance|
BBC Red Button 1|1464024300|The Super League Show|||0|0|Rugby League - Domestic|Tanya Arnold introduces action from the latest round of Super League matches, which saw every fixture take place at St James' Park in Newcastle on `Magic Weekend'.(n)
BBC Red Button 1|1464029700|EastEnders: Bobby: The Story So Far|||0|0|Soap,Melodrama|
BBC Radio 1|1463875200|DJ Target|||0|0||The home of new talent.(r)
BBC Radio 1|1463886000|Diplo and Friends|||0|0||Dance music.(r)
BBC Radio 1|1463893200|Dev|||0|0||Music and chat for Sunday morning.(r)
BBC Radio 1|1463907600|The Matt Edmondson Show|||0|0||Music and chat.(r)
BBC Radio 1|1463918400|Alice Levine|||0|0||Music and chat.(r)
BBC Radio 1|1463929200|Cel Spellman|||0|0||Your essential guide to the week, with great new pop and best bits from Radio 1, CBBC and online. Plus, from 6, it's the Number 1's Show.(r)
BBC Radio 1|1463940000|Rock Show with Daniel P Carter|||0|0||The best in modern and classic rock, including a round-up of the latest stories.(r)
BBC Radio 1|1463950800|Phil Taggart|||0|0||Music and chat.(r)
BBC Radio 1|1463961600|Monki|||0|0||Music from all corners of the club, featuring house and grime.(r)
BBC Radio 1|1463972400|Adele Roberts|||0|0||A selection of new and old music, as well as gossip and entertainment news.(r)
BBC Radio 1|1463981400|The Radio 1 Breakfast Show with Nick Grimshaw|||0|0||Craig David and Dan from Bastille take over the Radio 1 Breakfast Show in the run-up to the Big Weekend.(r)
BBC Radio 1|1463994000|Clara Amfo|||0|0||With chat, interviews and music from the Live Lounge.(r)
BBC Radio 1|1464003900|Newsbeat|||0|0||Headlines from around the world.(r)
BBC Radio 1|1464004800|Scott Mills|||0|0||A rousing mix of music, chat, competitions and entertainment news.(r)
BBC Radio 1|1464015600|Greg James|||0|0||Music, chat, competitions and entertainment news. Includes Newsbeat at 5.45pm.(r)
BBC Radio 1|1464026400|Annie Mac|||0|0||Music and chat.(r)
BBC Radio 1|1464033600|Radio 1's Playlists|||0|0||A guest selects music for their perfect playlists.(r)
BBC Radio 1|1464037200|Huw Stephens|||0|0||The DJ presents the best in new, unsigned and underground music from the UK and beyond.(r)
BBC Radio 1|1464048000|Friction|||0|0||Drum 'n' bass.(n)
BBC Radio 1|1464058800|Adele Roberts|||0|0||A selection of new and old music, as well as gossip and entertainment news.(n)
BBC Radio 1|1464067800|The Radio 1 Breakfast Show with Nick Grimshaw|||0|0||Jess Glynne and Ryan from OneRepublic take over the Radio 1 Breakfast Show. Plus, an appearance from Dominic Cooper.(n)
BBC Radio 1|1464080400|Clara Amfo|||0|0||With chat, interviews and music from the Live Lounge.(n)
BBC Radio 1|1464090300|Newsbeat|||0|0||Headlines from around the world.(n)
BBC Radio 1|1464091200|Scott Mills|||0|0||A rousing mix of music, chat, competitions and entertainment news.(n)
BBC Radio 1|1464102000|Greg James|||0|0||Music, chat, competitions and entertainment news. Includes Newsbeat at 5.45pm.(n)
BBC Radio 1|1464112800|Annie Mac|||0|0||Music and chat.(n)
BBC Radio 1|1464120000|Radio 1's Stories|||0|0||Clara Amfo and Dr Hannah Fry use numbers to explore the singer's career.(n)
BBC Radio 1|1464123600|Huw Stephens|||0|0||The DJ presents the best in new, unsigned and underground music from the UK and beyond.(n)
BBC Radio 2|1463882400|Bob Harris Sunday|||0|0||The host introduces a session performance by folk outfit Applewood Road, featuring Emily Barker, Amber Rubarth and Amy Speace.(r)
BBC Radio 2|1463893200|The Sunday Hour|||0|0||Diane Louise Jordan explores and celebrates diversity in the context of Trinity Sunday. She introduces readings and prayers as well as listeners' requests and dedications.(r)
BBC Radio 2|1463896800|Good Morning Sunday with Clare Balding|||0|0||The host presents a show focusing on ethical and religious issues, with contributions by her faith guest the Very Rev David Monteith, Dean of Leicester.(r)
BBC Radio 2|1463904000|Steve Wright's Sunday Love Songs|||0|0||A blend of love songs, dedications and real-life stories for romantics everywhere.(r)
BBC Radio 2|1463911200|The Michael Ball Show|||0|0||The broadcaster presents his regular Sunday lunchtime mix of music and chat, with TV and film previews, and a look at the day's papers.(r)
BBC Radio 2|1463918400|Elaine Paige on Sunday|||0|0||Musical theatre star Elaine Paige celebrates the sounds of Broadway, Hollywood and the West End.(r)
BBC Radio 2|1463925600|Johnnie Walker's Sounds of the 70s|||0|0||Johnnie is joined in conversation by Grammy Award-winning singer Rita Coolidge, and presents the usual mix of hits, album tracks and obscure tunes from the decade.(r)
BBC Radio 2|1463932800|Paul O'Grady|||0|0||The broadcaster introduces Triples featuring Frankie Goes to Hollywood and The Hollies. Plus, another hard-to-find old TV theme.(r)
BBC Radio 2|1463940000|Claudia on Sunday|||0|0||Two hours of requests, soundtrack choices and listener dedications. Plus the Great Sunday Songbook and Sunday Soak.(r)
BBC Radio 2|1463947200|Clare Teal|||0|0||The jazz singer presents a nostalgic review of the age of swing, featuring music by the big bands of Britain and America, from Benny Goodman to Quincy Jones.(r)
BBC Radio 2|1463954400|Moira Stuart|||0|0||The veteran broadcaster selects easy-listening tracks, including hits by Dianne Reeves, Melody Gardot, Jimmy Witherspoon and Matt Monro. Plus, an encounter between pianist Chick Corea and vibraphonist Gary Burton.(r)
BBC Radio 2|1463958000|After Midnight|||0|0||Music and chat with Janice Long, including Pause for Thought at 12.15am and 2.30am.(r)
BBC Radio 2|1463968800|Sounds of the 60s|||0|0||Brian Matthew presents chart hits and rarities from the early years of pop, including Marlena Shaw's Wade in the Water, and tracks from The Move's first album.(r)
BBC Radio 2|1463976000|Vanessa Feltz|||0|0||Early-morning music and chat. Including Pause for Thought at 5.45.(r)
BBC Radio 2|1463981400|Chris Evans|||0|0||Fun-packed show featuring music, entertainment and celebrity guests dropping by for a chat. Plus, sport and regular travel updates. Including at 9.15 Pause for Thought.(r)
BBC Radio 2|1463992200|Ken Bruce|||0|0||Jazz-infused pop singer Mari Wilson, known as the Neasden Queen of Soul, joins Ken to select her Tracks of My Years this week, beginning with hits by The Hollies and Abba.(r)
BBC Radio 2|1464001200|Jeremy Vine|||0|0||The broadcaster presents current-affairs chat live from the village of Dent in Cumbria, where asks residents whether they believe their community would benefit from a `Brexit'.(r)
BBC Radio 2|1464008400|Steve Wright in the Afternoon|||0|0||Music and chat, including Factoids, Non-Stop Oldies and the latest entertainment news.(r)
BBC Radio 2|1464019200|Simon Mayo|||0|0||Music, guests and discussion, with sports updates, the daily money feature and travel news.(r)
BBC Radio 2|1464026400|Paul Jones|||0|0||A selection of classic R&B tracks, including music by Young Jessie and Doug Sahm. Plus, a tribute to blues-rock guitarist and singer Lonnie Mack, who died on April 21.(r)
BBC Radio 2|1464030000|Jo Whiley|||0|0||The host reviews new releases by Eric Clapton, Catfish & the Bottlemen and Richard Ashcroft. Plus, the usual selection of Taxi Service dedications.(r)
BBC Radio 2|1464037200|Sounds of the 50s with Leo Green|||0|0||The musician and broadcaster celebrates musical gems from the 1950s, including tracks from a wide range of genres, from rock `n' roll to soul and swing.(r)
BBC Radio 2|1464040800|Jools Holland|||0|0||Songwriter, musician, producer and conductor Mike Batt joins Jools and his Rhythm and Blues Orchestra to chat about his career, and introduce some of his favourite music.(r)
BBC Radio 2|1464044400|After Midnight|||0|0||Music and chat with Janice Long, including Pause for Thought at 12.15am and 2.30am.(n)
BBC Radio 2|1464055200|Johnnie Walker's Sounds of the 70s|||0|0||Johnnie is joined in conversation by Grammy Award-winning singer Rita Coolidge, and presents the usual mix of hits, album tracks and obscure tunes from the decade.(n)
BBC Radio 2|1464062400|Vanessa Feltz|||0|0||Early-morning music and chat. Including Pause for Thought at 5.45.(n)
BBC Radio 2|1464067800|Chris Evans|||0|0||Music, features and celebrity guests. With sport and regular travel updates. Including Pause for Thought at 9.15.(n)
BBC Radio 2|1464078600|Ken Bruce|||0|0||The Neasden Queen of Soul Mari Wilson introduces her next two Tracks of My Years, highlighting music by Carole King and Mott the Hoople.(n)
BBC Radio 2|1464087600|Jeremy Vine|||0|0||The broadcaster's nationwide tour continues as he reaches Huddersfield, West Yorkshire, where he asks residents whether they believe their town would benefit from a `Brexit'.(n)
BBC Radio 2|1464094800|Steve Wright in the Afternoon|||0|0||New and vintage music, quirky facts and entertainment news.(n)
BBC Radio 2|1464105600|Simon Mayo|||0|0||Kenneth Branagh joins Simon to discuss the return of the English-language interpretation of Swedish detective drama Wallander, which premiered on BBC Four on Sunday.(n)
BBC Radio 2|1464112800|Jamie Cullum|||0|0||The pianist and songwriter presents interviews with Herbie Hancock, Chick Corea, Robert Glasper and others recorded at the White House in Washington, DC on International Jazz Day.(n)
BBC Radio 2|1464116400|Jo Whiley|||0|0||A mix of new music and classic tracks, with guests dropping in to the studio to chat.(n)
BBC Radio 2|1464123600|Paper Cuts|||0|0||Kate Thornton invites more celebrity guests to revisit landmark events from their careers via print headlines, beginning with broadcaster Gloria Hunniford.(n)
BBC Radio 2|1464127200|Nigel Ogden: The Organist Entertains|||0|0||Organs in a variety of grand settings including Liverpool's Anglican Cathedral, Hull City Hall and Trono Church in Sweden, featuring Graham Barber, David Poulter and Carlo Curley.(n)
BBC Radio 2|1464129000|Listen to the Band|||0|0||Frank Renton introduces more music from the Gala Concert at the European Brass Band Championships in Lille, featuring The Black Dyke Band, and the European Youth Brass Band.(n)
BBC Radio 3|1463871600|Geoffrey Smith's Jazz|||0|0||Geoffrey Smith revisits the music of Dexter Gordon and Wardell Gray, who were renowned as `bebop's tenor kings' famed for their saxophone duels. Geoffrey recalls those thrilling encounters, and their later individual careers.(r)
BBC Radio 3|1463875200|Through the Night|||0|0||With Catriona Young. Haydn: Sinfonia concertante in B flat, H1 105 for oboe, bassoon, violin, cello and orchestra. Hélène Devilleneuve (oboe), Jean-François Duquesnoy (bassoon), Hélène Collerette (violin), Daniel Racolt (cello), Radio France Philharmonic Orchestra, conducted by Ton Koopman. 1.23 Bach: Concerto in C minor for oboe, violin and strings, BWV1060R (reconstr Schneider). 1.36 Handel: Concerto a due cori No 3 in F, HWV334. 1.52 Daniel-Lesur: Le Cantique des colonnes. 2.05 Messiaen: Quatuor pour la fin du temps for clarinet, piano, violin and cello. 2.54 Melartin: Lohdutus (Consolation). 3.01 Schubert: Six Moments musicaux for piano, D780. 3.30 Beethoven: Symphony No 1 in C, Op 21. 3.59 Telemann: Affetuoso and aria: Wandelt in der Liebe, gleich wie Christus uns geliebt! 4.06 Kalnins: Ballad for cello and piano. 4.13 Jommelli: Sonata in D. 4.23 Liszt: La Campanella. 4.29 Mozart: Duet: Fra gli amplessi (Così fan tutti). 4.35 Auber: Overture to Marco Spada. 4.46 Vivaldi: Concerto for bassoon and orchestra in A minor, RV497. 5.01 Ruth Watson Henderson: Come Holy Spirit for SATB with organ accompaniment. 5.06 Förster: Jesu dulcis memoria. 5.13 Chopin: Two Nocturnes for piano, Op 27: No 1 in C sharp minor; No 2 in D flat. 5.26 Salmenhaara: Adagietto for Orchestra (1981). 5.32 Britten: A Charm of lullabies for mezzo-soprano and piano, Op 41. 5.44 Ibert:Trio for violin, cello and harp. 5.59 Grieg: Peer Gynt: Suite No 1, Op 46. 6.24 Meulemans: Five Piano Pieces: Als de beke zingt (When the brook is chanting); Menuet; Mazurka triste; Wals; Lentewandeling (Vernal wanderings). 6.43 Bach: Quartet for flute, viola and continuo in D, Les Adieux, Andreas Staier (fortepiano), Wilbert Hazelzet (flute), Hajo Bäß (viola).(r)
BBC Radio 3|1463896800|Breakfast|||0|0||Music, news and the occasional surprise, presented by Elizabeth Alker. Including 7.00, 8.00 News.(r)
BBC Radio 3|1463904000|News|||0|0||
BBC Radio 3|1463904180|Sunday Morning with James Jolly|||0|0||Prompted by this week's Building A Library selection, Handel's Alcina, Jonathan Swain looks at how other composers have depicted sorcery and magic, from Handel's contemporary Caldara to Ligeti, by way of Dukas and Janácek. The young artist spotlight is on harpsichordist Maxim Emelyanychev, and the British masterpiece of the week is Elgar's Introduction and Allegro for Strings, Op 47.(r)
BBC Radio 3|1463914800|Private Passions|||0|0||Jane Goodall was only twenty-four when in she went to live among the chimpanzees of Gombe National Park in Tanzania, and she went on to spend more than 55 years there. She has done more than anyone else to transform our understanding of chimpanzees - and beyond that, her work has raised questions about how we treat these highly intelligent primates, and indeed about the rights of all animals. Now in her early eighties, she's on an extraordinary mission travelling round the world to protect chimpanzees from extinction. During a rare stay in Britain, Jane Goodall talks to Michael Berkeley about her life and ground-breaking discoveries. She reveals that the chimpanzees she lived with also had a darker side, and were sometimes violent, stamping on her. She remembers difficult times after the kidnapping of some of her workers, and the death of her second husband and how music sustained her, and transformed her view of the world. Music choices include Beethoven, Bach, Schubert, Mendelssohn's Violin Concerto and Richard Burton reading the Dylan Thomas classic Under Milk Wood. She also introduces some very excited chimpanzee speech, and speculates about what kind of music chimpanzees enjoy.(r)
BBC Radio 3|1463918400|News|||0|0||
BBC Radio 3|1463918520|Radio 3 Lunchtime Concert|||0|0||The Jerusalem Quartet performs quartets by Beethoven and Bartok from Wigmore Hall, London. Beethoven builds the elaborate first and second movements of his Op 18 No 2, from a simple melodic idea, while Bartok prefaces his String Quartet No 6 with the same melancholy theme and uses it as the basis of the work as introspective finale. Beethoven: String Quartet in G, Op 18, No 2. Bartok: String Quartet, No 6.(r)
BBC Radio 3|1463922000|The Early Music Show|||0|0||Hannah French presents highlights of a concert given by the Flanders Recorder Quartet at The Frick Collection in New York, including music by JS Bach, Hugh Ashton, Tielman Susato and Joseph de Boismortier. Hannah also talks to artistic director Joyce Bodig about the museum's long-standing series of chamber music concerts and talks to chief curator Xavier Salomon about some of the works of art in the collection.(r)
BBC Radio 3|1463925600|Choral Evensong|||0|0||Live from Tewkesbury Abbey and sung by the Abbey's Schola Cantorum. Introit: Gracious Spirit, Holy Ghost (Sebastian Forbes). Responses: Richard Shephard. Psalms 93, 94 (Bell, Deffell (after Cherubini), Peterson). Office Hymn: Breathe on me, Breath of God (Carlisle). First Lesson: Genesis 15. Canticles: Westminster Service (Howells). Second Lesson: Romans 4 vv.1-8. Anthem: Dum complerentur (Palestrina). Final Hymn: Come down, O Love divine (Down Ampney). Organ Voluntary: Tongues of Fire (Arthur Wills) Director: Simon Bell. Organist: Carleton Etherington.(r)
BBC Radio 3|1463929200|The Choir|||0|0||Sara Mohr-Pietsch meets a group of singers who also have a love of gardening at the Chelsea Flower Show. Plus, a look ahead to Harrogate-based barbershop festival Sing 2016.(r)
BBC Radio 3|1463932800|The Listening Service|||0|0||The Listening Service - an odyssey through the musical universe with Tom Service. Join him on a journey of imagination and insight, exploring how music works. Today - What's all that that Noise? Tom investigates - when is noise just noise, and when is it music? is it just sound in the wrong place? Tom finds that, though we resent noises in the concert hall, music needs some noise in it to give it character. He also investigates the contemporary genre of Noise Music at an avant garde club. He considers noise in our daily lives, and talks to Emily Cockayne, author of Hubbub: Filth Noise & Stench in England 1600-1770; and to David Hendy, author of Noise: a Human History. We can't avoid noise, so can we learn to love it?.(r)
BBC Radio 3|1463934600|Words and Music|||0|0||The baobab tree is one of the most recognisable species in Africa. In many places, the enduring giant trees are a symbol of community, a place of gathering, and a location to exchange stories. Storytelling has played a fundamental role in communities across Africa for centuries, with the oral traditions of myths and legends handed down through generations. In modern times poets and writers have often focussed on the effects of colonialism, recent conflicts, and questions of identity. Combining these demonstrates the richness of African literature and the issues facing different nations today. Including music from Africa and beyond.(r)
BBC Radio 3|1463939100|Sunday Feature|||0|0||Michael Goldfarb tells the story of Dutch philosopher Benedict Spinoza, who 350 years ago, asked Who is God? and what role should religion play in government. In the middle of 17th century Europe religion and politics were inseparable and the result was bloodshed everywhere. Then a Dutch Jew, Benedict Spinoza, wrote a book that challenged this idea of government. His argument: get priests and clergy out of politics. People should not be ruled by monarchs who claimed they were anointed by God. Let there be democracy, where reason and intellect guide the state. You can guess how this argument was received. Spinoza was called 'the renegade Jew from Hell.' Michael Goldfarb tells the story of this God Intoxicated Man and the world in which he lived - the Golden Age of the Dutch Republic - and how he has become the philosopher with new relevance for our times. Atheist, pantheist, heretic, or none of those things; man of science and moral philosopher, Spinoza's conception of the universe has influenced scientists, playwrights, novelists, poets and musicians. Using Spinoza's own words, interviews with philosophers and music inspired by his thoughts, Goldfarb tells the story of the man of whom it was said, 'Christ was sent to redeem man. Spinoza was born for a far greater purpose. He was born to redeem God.'.(r)
BBC Radio 3|1463941800|Radio 3 in Concert|||0|0||Nikolaus Harnoncourt conducts Concentus Musicus in two Viennese masterpieces. The Austrian conductor is heard here in two of his last concerts where his typically inspirational performances with his own period instrument orchestra are a reminder of why he is seen as one of the most influential musicians of the past half century. Presented by Ian Skelly. Haydn: Mass No. 10 in C, Hob. XXII:9 ('Missa in Tempore Belli') ('Paukenmesse'). Sylvia Schwartz (soprano), Elisabeth von Magnus (mezzo-soprano), Daniel Johannsen (tenor), Ruben Drole (bass), Arnold Schoenberg Choir, Concentus Musicus, Vienna, conductor Nikolaus Harnoncourt, rec. Parish Church, Stainz - Styriarte Festival - 12.07.15. Beethoven: Symphony No. 5 in C minor, op. 67. Concentus Musicus, Vienna, conductor Nikolaus Harnoncourt, rec. Musikverein, Vienna - 10.05.15.(r)
BBC Radio 3|1463947200|Drama on 3|||0|0||What happened to Jessica, Shylock's daughter in The Merchant of Venice? In the original Shakespeare, Jessica is a minor but fascinating character, Shylock's only daughter, who leaves him to convert to Christianity and marry Lorenzo. We are left rather uncertain about how that marriage is going to work out. It's also implicit that the conversion isn't going to be easy on either party. The Wolf in the Water by Naomi Alderman is an imaginative response to The Merchant of Venice, in which we meet an older Jessica in 1615, secretly still practising her Jewish faith in a turbulent Venice that is increasingly hostile to Jews. A murder, twenty innocent Jews facing death - Jessica becomes embroiled in a mystery that challenges her apparently settled life and reconnects her with her identity. The year may be 1615, but the themes are universal and relevant. What drives one group to persecute another? What shameful deeds are done by those to whom we entrust our money? Can we ever be cosmopolitans - citizens of all nations and none - or will our ethnicity, our religion, even the ineradicable traces of God, always draw us back, perhaps to doom ourselves? Naomi Alderman is an award-winning writer, writing her first BBC Radio 3 drama commission, after establishing herself at the cutting edge of new fiction and audio gaming. Part of the BBC's Shakespeare Festival but also marking the 500th anniversary of the establishment of the Venice ghetto.(r)
BBC Radio 3|1463952600|Early Music Late|||0|0||Elin Manahan Thomas presents a performance of Handel's Water Music performed by the Akademie fur Alte Musik Berlin at the Amsterdam Concertgebouw earlier this year. Handel: Water Music, HWV 348-350. Akademie fur Alter Musik Berlin, Georg Kallweit (director/violin).(r)
BBC Radio 3|1463956200|Britten in Venice|||0|0||Britten's String Quartet No 3, performed by the Amadeus Quartet and his Suite: Death in Venice, arranged and conducted by Steuart Bedford, both pieces inspired by the great city in which he spent much time during his latter years.(r)
BBC Radio 3|1463959800|Through the Night|||0|0||With Catriona Young. 12.31Schubert: Symphony no.4 in C minor, D.417 'Tragic'. 12.58 Bruckner: Mass no.3 in F minor for soloists, chorus, orchestra and organ. 2.01 Sibelius: Symphony no.7 (Op.105) in C major. 2.22 Liszt: Sonetto 123 di Petrarca (S.158 No.3): Io vidi in terra angelici costumi. 2.31 Beethoven:Trio for strings (Op.9`1) in G major. 3.00 Grieg:Haugtussa - song cycle. 3.27 Borodin: Polovtsian dances from 'Prince Igor'. 3.38 Chopin: Three Mazurkas (Op.59). 3.49 Pandolfi Mealli: Sonata in E minor Op.4`1 (La Bernabea) for violin and continuo. 3.55 JS Bach: 6 Chorales from the Schemelli Collection: Gott, wie gross ist deine Güte (BWV.462); Dich bet' ich an, mein höchster Gott (BWV.449); Dir, dir, Jehova, will ich singen (BWV.452); O liebe Seele, zieh' die Sinnen (BWV.494); Vergiss mein nicht, mein allerliester Gott (BWV.505); Ich halte treulich still und liebe meinen Gott (BWV.466). 4.08 Vivaldi: Concerto da Camera in C major (RV.88). 4.15 Chaminade: Concertino Op.107. 4.24 Dvorák: Slavonic Dance No.10 in E minor (Op.72 No.2) (Starodávny). 4.31 Mozart: Kirchen-Sonate in B flat (K. 212) for 2 violins, double bass and organ. 4.36 Field: Andante inédit in E flat major for piano. 4.44 Haydn: Trio in E flat major H.15.30 for keyboard and strings. 5.02 Bach: Siehe, wie fein und lieblich ist es - vocal concerto for 2 tenors, bass and instruments. 5.09 Boccherini: La Musica Notturna delle strade di Madrid Quintet No 6, Op 30 (G.324). 5.22 Guerau: Mariona from 'Poema Harmonico'. 5.28 Debussy: Iberia - from Images for Orchestra. 5.49 Rachmaninov: Suite for 2 pianos in G minor (Op.5) (Fantasie-Tableaux). 6.15 Locatelli: Violin Concerto in E flat (Op.7 No.6), 'Il Pianto d?Arianna'.(r)
BBC Radio 3|1463981400|Breakfast|||0|0||Music, news and the occasional surprise, presented by Petroc Trelawny. Including 7.00, 8.00 News. 7.30, 8.30 News Headlines.(r)
BBC Radio 3|1463990400|Essential Classics|||0|0||With Rob Cowan. 9.00 My favourite... Handel Concerti Grossi Op. 6. Rob shares his favourite baroque masterpieces from Handel's 12 grand concertos, features performances of them by the Academy of Ancient Music, Concentus Musicus Wien, Il Giardino Armonico and the Boyd Neel Orchestra. 9.30 The daily musical challenge is to name the film or TV programme that featured a certain piece of classical music. 10.00 Rob's guest is author Malorie Blackman, who has written more than 60 books for children and young readers and was the Children's Laureate from 2013 to 2015. Malorie shares a selection of her favourite classical music, including works by the 19th-century composer Samuel Coleridge Taylor, and Florence Price, the first African-American woman to have a composition performed by a major symphony orchestra.10:30 Music in Time. The focus is on the Medieval period and the great chanson composer Clément Janequin, whose song La chant des oiseaux imitates birdsong. 11.00 The Artist of the Week is the Suk Trio, with recordings including Mendelssohn's Piano Trio in D Minor Op. 49, Dvorak's Piano Trio No.3 in F minor, Op.65 and Brahms's Piano Trio No.1 in B major, Op.8. Mendelssohn: Piano Trio in D minor, Op.49. Suk Trio.(r)
BBC Radio 3|1464001200|Composer of the Week: Clara Schumann and Her Circle|||0|0||Donald Macleod explores the lives and music of Clara Schumann and the composers and musicians whose circles she moved in, beginning with Chopin. Clara was 13 when she first encountered Chopin in the early months of 1832 during a promotional visit to Paris and she was in the audience for his astonishing first public Parisian recital, at the Salle Pleyel. She had already learnt one of his works, and his music would be a mainstay of her concert repertoire for the next six decades. The respect was clearly mutual as when Chopin visited Clara in Leipzig a few years later, he was impressed enough to take several of her pieces away with him. C Schumann: 4 Polonaises, Op 1 (No 2 in C). Suzanne Grutzmann (piano). Chopin: Variations on Mozart's Là ci darem la mano, Op 2. Garrick Ohlsson (piano), Warsaw Philharmonic Orchestra, conductor Kazimierz Kord. C Schumann: Soirées musicales, Op 6 (No 4, Ballade in D minor); 4 Pièces caracteristiques, Op 5 (No 4, Scène fantastique (Le ballet des Revenants)). Suzanne Grutzmann (piano). Chopin: Cello Sonata in G minor, Op 65 (3rd mvt, Largo). Mischa Maisky (cello), Martha Argerich (piano). C Schumann: Piano Concerto in A minor, Op 7 (3rd mvt, Finale. Allegro non troppo). Lucy Parham (piano), BBC Concert Orchestra, conductor Barry Wordsworth.
BBC Radio 3|1464004800|News|||0|0||
BBC Radio 3|1464004920|Radio 3 Lunchtime Concert|||0|0||Sara Mohr-Pietsch presents from London's Wigmore Hall as violinist Pekka Kuusisto and cellist Nicolas Altstaedt perform arrangements of Two-part inventions by Bach, duos by contemporary German composer Jörg Widmann and Ravel's Sonata, a classic for this combination of instruments. Bach: Two-part Inventions (selection). Jörg Widmann: 24 Duos (selection). Ravel: Sonata for violin and cello. Pekka Kuusisto (violin), Nicolas Altstaedt (cello).(r)
BBC Radio 3|1464008400|Afternoon on 3|||0|0||Verity Sharp presents the first of a week of programmes featuring the BBC National Orchestra of Wales, including an archive performance from Leningrad in 1988. 2.00 Walton: Portsmouth Point. BBC National Orchestra of Wales, conductor Rumon Gamba. 2.05 Tchaikovsky: Romeo and Juliet - fantasy overture. Conductor Thomas Sondergard. 2.25 Rachmaninov: Piano Concerto no. 2 in c minor op. 18. Freddy Kempf (piano), conductor Thomas Sondergard. 3.05 Prokofiev: Romeo and Juliet [sel. Sondergard]. Conductor Thomas Sondergard. 3.55 Strauss: Don Juan. Conductor Tadaaki Otaka. 4.15 Mussorgsky: Night on the Bare Mountain. Conductor Grant Llewellyn.(r)
BBC Radio 3|1464017400|In Tune|||0|0||Sean Rafferty is joined by guitarist Sean Shibe, who performs live ahead of his appearance at Bath International Music Festival. Including 5.00, 6.00 News.(r)
BBC Radio 3|1464024600|Composer of the Week: Clara Schumann and Her Circle|||0|0||Donald Macleod explores the lives and music of Clara Schumann and the composers and musicians whose circles she moved in, beginning with Chopin. Clara was 13 when she first encountered Chopin in the early months of 1832 during a promotional visit to Paris and she was in the audience for his astonishing first public Parisian recital, at the Salle Pleyel. She had already learnt one of his works, and his music would be a mainstay of her concert repertoire for the next six decades. The respect was clearly mutual as when Chopin visited Clara in Leipzig a few years later, he was impressed enough to take several of her pieces away with him. C Schumann: 4 Polonaises, Op 1 (No 2 in C). Suzanne Grutzmann (piano). Chopin: Variations on Mozart's Là ci darem la mano, Op 2. Garrick Ohlsson (piano), Warsaw Philharmonic Orchestra, conductor Kazimierz Kord. C Schumann: Soirées musicales, Op 6 (No 4, Ballade in D minor); 4 Pièces caracteristiques, Op 5 (No 4, Scène fantastique (Le ballet des Revenants)). Suzanne Grutzmann (piano). Chopin: Cello Sonata in G minor, Op 65 (3rd mvt, Largo). Mischa Maisky (cello), Martha Argerich (piano). C Schumann: Piano Concerto in A minor, Op 7 (3rd mvt, Finale. Allegro non troppo). Lucy Parham (piano), BBC Concert Orchestra, conductor Barry Wordsworth.
BBC Radio 3|1464028200|Radio 3 in Concert|||0|0||Jamie MacDougall presents a concert from Glasgow's City Halls in which Donald Runnicles conducts the BBC SSO in Mahler's Symphony No 1 and soloist Denis Kozhukhin joins them for Brahms' Piano Concerto No 2. There has never been a first symphony to match Mahler's, from the glistening stillness of its visionary opening to its final, epic ascent from the inferno to paradise. It is a suitably joyous ending to the orchestra's 80th anniversary season and to a concert that begins with the poetry and warmth of Brahms's expansive Second Piano Concerto: a Romantic master at his big-hearted best, and a glowing conclusion to Denis Kozhukhin's BBC SSO Brahms cycle. Brahms: Piano Concerto No 2. 8.20 Interval. 8.40 Mahler: Symphony No 1. BBC Scottish Symphony Orchestra, Donald Runnicles (conductor) Denis Kozhukhin (piano).(r)
BBC Radio 3|1464037200|Music Matters|||0|0||Tom Service with a portrait of the Romanian composer George Enescu, as his masterpiece opera Oedipe is staged for the first time at the Royal Opera House in London. Among the contributors are Professor Erik Levi, expert on music of the 20th-Century; the Romanian violinist Remus Azoitei, and the American conductor Lawrence Foster, former director of the Enescu Festival in Bucharest. Also, Tom interviews pianist Steven Osborne on the parallels and differences between George Crumb and Morton Feldman, two American modernist composers obsessed with new sounds and textures in music. Also, the composer Philip Venables on his opera 4.48 Psychosis, based on the iconic play by Sarah Kane exploring depression - the first ever adaptation of her work on stage, to be premiered this month at the Lyric Hammersmith in London.(r)
BBC Radio 3|1464039900|The Essay|||0|0||Prominent people in a particular line of work read and reflect on the writings of an illustrious person who plied the same trade. In the first edition, teacher Francis Gilbert reads Jean-Jacques Rousseau's Emile's and assesses whether this template for a perfect education has a place and an influence on today's curriculum.(r)
BBC Radio 3|1464040800|Jazz Now|||0|0||Soweto Kinch presents the UK premiere of Julian Arguelles' suite of South African-inspired music with Steve Arguelles, Django Bates and Frankfurt Radio Big Band recorded at the Cheltenham Jazz Festival.(r)
BBC Radio 3|1464046200|Through the Night|||0|0||With Catriona Young. 12. 31 Tchaikovsky: Jurists' March in D. 12.37 Scriabin: Piano Concerto No.1 in F sharp minor, Op.20. 1.05 Scriabin: Piano Sonata No.4 in F sharp major, Op.30. 1.13 Glazunov: The Seasons - ballet in one act, Op.67. 1:51Vladigerov: Elegie d'automne - from 3 pieces pour piano (Op.15). 1.58 Pipkov: Nani mi nani, Damiancho. 2.03 Kandov: Trio-concerto for Harp, Flute, Cello and String Orchestra. 2.26 Kutev: Dragana and the Nightingale. 2.31Vladigerov: Divertimento for chamber orchestra. 2.47 Prokofiev, arr. Prokofiev & David Oistrakh: Sonata for violin and piano No.2 (Op.94bis) in D major. 3.13 Delibes: Entracte from 'Lakmé'. 3.17 Delibes: Couplets de Nilacantha de l'acte II de l'opera 'Lakmé'. 3:21 Strauss: An einsamer Quelle from Stimmungsbilder (Op.9 No.2); Intermezzo from Stimmungsbilder (Op.9 No.3). 3.30 Hristov: Heruvimska pesen no.4 (Cherubic Song). 3.37 JS Bach & Gounod: Ave Maria (arr. for trumpet and organ by Blagoj Angelovski). 3.46 Busoni: Concertino for clarinet and small orchestra (Op.48) in B flat major. 3:58 Dvorák: Romance (Op.11) in F minor vers. for violin and piano. 4.10 Dinev: Milost mira No.6 (A Mercy of Peace No.6). 4.15 JS Bach: Concerto for oboe d'amore and string orchestra No.4 (BWV.1055) in A major. 4.31 Infante:Three Andalucian Dances. 4.46 Anonymous:Folias de Espana. 4.53 Granados, arr. Chris Paul Harman: La Maja y el Ruiseñor - from Goyescas. 5.00 Handel: Spirit Music (Nos.1 to 4) - from Alcina. 5.07 Schubert: Quartettsatz for strings in C minor (D.703). 5.17 Brahms: Marienlieder (Op.22). 5.35 Bach: Sonata for violin and harpsichord in B minor (H.512). 5.53 Crusell: Concertino for bassoon and orchestra in B flat major. 612 Liszt: Liebestraume (S.541) no.3 in A flat major. 6:18 Janácek: Pohádka for cello and piano.(n)
BBC Radio 3|1464067800|Breakfast|||0|0||Petroc Trelawny presents Radio 3's classical breakfast show, featuring listener requests. Including 7.00, 8.00 News. 7.30, 8.30 News Headlines.(n)
BBC Radio 3|1464076800|Essential Classics|||0|0||With Rob Cowan. 9.00 My favourite Handel Concerti Grossi, Op 6. Rob shares his favourite Baroque masterpieces from Handel's Twelve Grand Concertos. The line-up features performances of these energetic concertos by the Academy of Ancient Music directed by Andrew Manze, Concentus Musicus Wien and Nikolaus Harnoncourt, Il Giardino Armonico under Giovanni Antonini, and Thurston Dart conducting the Boyd Neel Orchestra. 9.30 A musical challenge to identify a piece of music played backwards. 10.00 Rob's guest is author Malorie Blackman, who shares a selection of her favourite classical music. 10.30 Music in Time: Modern. Rob explores the Modern period with Bartok's Music for Strings, Percussion and Celesta, a score that reignited a fascination with spatially separated musicians. 11.00 Rob's Artist of the Week is the Suk Trio. Throughout the week Rob delves into the archives of this internationally renowned piano trio, sharing recordings including Mendelssohn's Piano Trio in D minor, Op 49, Dvorak's Piano Trio No 3 in F minor, Op 65 and Brahms's Piano Trio No 1 in B major, Op 8. Dvorak: Piano Trio No 3 in F minor, Op 65. Suk Trio.(n)
BBC Radio 3|1464087600|Composer of the Week: Clara Schumann and Her Circle|||0|0||Donald Macleod explores the lives and music of Clara Schumann and the extraordinary circle of composers and musicians she moved in. Much of Robert Schumann's music is a love-letter to Clara, translating key events in their relationship into sound - and from the start, Clara became its principal advocate and most authoritative interpreter. Clara Schumann: Soirées musicales, Op 6 (No 1, Toccatina in A minor). Jozef de Beenhouwer (piano). Soirées musicales, Op 6 (No 2, Notturno). Konstanze Eickhorst (piano). Robert Schumann: Novelletten, Op 21 (No 8, Sehr lebhaft (Stimme aus der Ferne)). Eric le Sage (piano). Clara Schumann: Am Strande; Warum willst du andre fragen, Op 12 No 11; Liebst du um Schönheit, Op 12 No 4; Er ist gekommen, Op 12 No 2. Christina Högman (soprano), Roland Pöntinen (piano). Robert Schumann: Six Etudes pour le pianoforte d'après les caprices de Paganini, Op 3 (No 1 in A minor; No 2 in E). Mariya Kim (piano). Clara Schumann: Variations on a Theme of Robert Schumann, Op 20. Jozef de Beenhouwer (piano).(n)
BBC Radio 3|1464091200|News|||0|0||
BBC Radio 3|1464091320|Radio 3 Lunchtime Concert|||0|0||Hannah French presents chamber music by Purcell, Haydn and Beethoven from the Frick Collection in New York. Cellist Nicolas Altstaedt and pianist Alexander Lonquich perform Beethoven's Seven Variations on 'Bei Männern welche Liebe fühlen', the Minetti Quartet plays Haydn's 'Sunrise' quartet, Op 76 No 4. Plus, there are songs by Purcell and Kate Bush from mezzo-soprano Anne-Sofie von Otter, with lutenist Thomas Dunford and keyboard player Jonathan Cohen.(n)
BBC Radio 3|1464094800|Afternoon on 3|||0|0||Verity Sharp presents music by the BBC National Orchestra of Wales, as baroque expert Rachel Podger directs from the violin in a Vivaldi concerto, and Damian Iorio makes his debut with the orchestra in music inspired by Italy. Recent Radio 3 New Generation Artist Olena Tokar returns to the orchestra with whom she sang at BBC Cardiff SInger of the World in 2013, with a setting of a poem by Shelley. Ansell: Plymouth Hoe. BBC National Orchestra of Wales, conductor Rumon Gamba. 2.10 Grace Williams: Sea Sketches, conductor Tadaaki Otaka. 2.30 Elgar: In the South (Alassio), conductor Thierry Fischer. 2.55 Vivaldi: Violin Concerto, Op 9 No 6, director Rachel Podger (violin). 3.05 Liszt: Legends, conductor Damian Iorio. 3.25 Respighi: Il Tramonto. Olena Tokar (soprano), conductor Damian Iorio. 4.00 Respighi: Church Windows, conductor Damian Iorio.(n)
BBC Radio 3|1464103800|In Tune|||0|0||Suzy Klein presents a programme to accompany the launch today of BBC Music Get Playing, which aims to boost amateur music-making around the country. Including 5.00, 6.00 News.(n)
BBC Radio 3|1464111000|Composer of the Week: Clara Schumann and Her Circle|||0|0||Donald Macleod explores the lives and music of Clara Schumann and the extraordinary circle of composers and musicians she moved in. Much of Robert Schumann's music is a love-letter to Clara, translating key events in their relationship into sound - and from the start, Clara became its principal advocate and most authoritative interpreter. Clara Schumann: Soirées musicales, Op 6 (No 1, Toccatina in A minor). Jozef de Beenhouwer (piano). Soirées musicales, Op 6 (No 2, Notturno). Konstanze Eickhorst (piano). Robert Schumann: Novelletten, Op 21 (No 8, Sehr lebhaft (Stimme aus der Ferne)). Eric le Sage (piano). Clara Schumann: Am Strande; Warum willst du andre fragen, Op 12 No 11; Liebst du um Schönheit, Op 12 No 4; Er ist gekommen, Op 12 No 2. Christina Högman (soprano), Roland Pöntinen (piano). Robert Schumann: Six Etudes pour le pianoforte d'après les caprices de Paganini, Op 3 (No 1 in A minor; No 2 in E). Mariya Kim (piano). Clara Schumann: Variations on a Theme of Robert Schumann, Op 20. Jozef de Beenhouwer (piano).(n)
BBC Radio 3|1464114600|Radio 3 in Concert|||0|0||The Royal Scottish National Orchestra, conducted by Peter Oundjian, perform a powerful Russian programme of Shostakovich's eighth symphony and Prokofiev's spirited second piano concerto, from Glasgow Royal Concert Hall. Presented by Tom Redmond. Nikolai Lugansky (piano), Royal Scottish National Orchestra, conductor Peter Oundjian. Prokofiev: Piano Concerto No 2. 8.05 Interval: Schubert: Four Impromptus, D935 performed by Nikolai Lugansky. 8.25 Shostakovich: Symphony No 8.(n)
BBC Radio 3|1464123600|Free Thinking|||0|0||Matthew Sweet talks to three photographers aged over 90 - Dorothy Bohm, Wolfgang Suschitzky and Neil Libbert - and to the inventor of the World Wide Web Tim Berners-Lee.(n)
BBC Radio 3|1464126300|The Essay|||0|0||Theatre critic Susannah Clapp explores Oscar Wilde's essay on criticism, finding that he was on the wrong side of anonymity arguments.(n)
BBC Radio 3|1464127200|Late Junction|||0|0||Nick Luscombe introduces music recorded live from the Late Junction stage at The Great Escape festival in Brighton. Plus, tracks by Portuguese-Angolan collective Throes + The Shine.(n)
BBC Radio 4 FM|1463871600|News and Weather|||0|0||
BBC Radio 4 FM|1463873400|Stories from Songwriters|||0|0||The first in a series of specially commissioned stories by songwriters, beginning with Sunset to Break Your Heart by Barb Jungr - a touching story that is set on the Shetland Islands. Read by Suranne Jones.(r)
BBC Radio 4 FM|1463874480|Shipping Forecast|||0|0||
BBC Radio 4 FM|1463875200|As BBC World Service|||0|0||
BBC Radio 4 FM|1463890800|Shipping Forecast|||0|0||
BBC Radio 4 FM|1463891400|News Briefing|||0|0||
BBC Radio 4 FM|1463892180|Bells on Sunday|||0|0||The morning bells from the Parish Church of St Thomas in Hazel Grove, Stockport, ringing Cambridge Surprise Major.(r)
BBC Radio 4 FM|1463892300|Profile|||0|0||Friends, adversaries, colleagues and confidants provide an insight into the personality and motivation of Ruth Davidson, leader of the Scottish Conservatives. Mark Coles presents.(r)
BBC Radio 4 FM|1463893200|News Headlines|||0|0||
BBC Radio 4 FM|1463893500|Something Understood|||0|0||Mark Tully examines deterrence, revealing how it often fails to work and can have harmful consequences by preventing people from pursuing other options.(r)
BBC Radio 4 FM|1463895300|Living World|||0|0||Archive programme in which Lionel Kelleway tracks down radio-tagged hedgehogs as they wake up from hibernation and enter into courtship rituals. Introduced by Chris Packham.(r)
BBC Radio 4 FM|1463896620|Weather|||0|0||
BBC Radio 4 FM|1463896800|News|||0|0||
BBC Radio 4 FM|1463897220|Sunday Papers|||0|0||Review of the latest news stories making the headlines.(r)
BBC Radio 4 FM|1463897400|Sunday|||0|0||Thomas Becket's relic; a new book giving voice to Transgender Christians and the World Humanitarian Summit, some of the stories in this week's programme.(r)
BBC Radio 4 FM|1463900100|Radio 4 Appeal|||0|0||Ian McEwan presents an appeal on behalf of SolarAid.(r)
BBC Radio 4 FM|1463900220|Weather|||0|0||
BBC Radio 4 FM|1463900400|News|||0|0||
BBC Radio 4 FM|1463900820|Sunday Papers|||0|0||Review of the latest news stories making the headlines.(r)
BBC Radio 4 FM|1463901000|Sunday Worship|||0|0||A Mass for Trinity Sunday live from St Anne's Cathedral, Leeds.(r)
BBC Radio 4 FM|1463903280|A Point of View|||0|0||Will Self questions whether the mind is stronger than the body, and what effect the ubiquity of psychiatrists and psychoanalysts plays in modern Britain.(r)
BBC Radio 4 FM|1463903880|Tweet of the Day|||0|0||Miranda Krestovnikoff presents the unusual chirring sound of the nightjar, a bird often heard calling on summer evenings.(r)
BBC Radio 4 FM|1463904000|Broadcasting House|||0|0||A discussion on the week's major headlines, presented by Paddy O'Connell.(r)
BBC Radio 4 FM|1463907600|The Archers|||0|0||Omnibus. Peggy makes a decision, and there is an awkward moment at the Bull.(r)
BBC Radio 4 FM|1463912100|Desert Island Discs|||0|0||Motown producer Berry Gordy talks to Kirsty Young and selects eight records to take to the mythical island.(r)
BBC Radio 4 FM|1463914800|News|||0|0||
BBC Radio 4 FM|1463915040|Just a Minute|||0|0||The comedy panel show returns for its 75th series, with Paul Merton, John Finnemore, Gyles Brandreth and Sheila Hancock joining host Nicholas Parsons as they try to speak on a given topic for 60 seconds without hesitation, repetition or deviation.(r)
BBC Radio 4 FM|1463916600|The Food Programme|||0|0||The first of two programmes in which author Diana Henry talks to Sheila Dillon about the writers who shaped her passion for food. With readings by Rebecca Ripley and Sam Woolf.(r)
BBC Radio 4 FM|1463918220|Weather|||0|0||
BBC Radio 4 FM|1463918400|The World This Weekend|||0|0||Global news and analysis, presented by Mark Mardell.(r)
BBC Radio 4 FM|1463920200|Jutland: The Battle that Won the War|||0|0||Lord Alan West explains why he believes Jutland was the most important First World War battle, a strategic victory that directly paved the way for allied victory.
BBC Radio 4 FM|1463922000|Gardeners' Question Time|||0|0||Eric Robson hosts a correspondence edition from Ness Botanic Gardens in The Wirral, where Christine Walkden, Bob Flowerdew and Pippa Greenwood answer listeners' queries.(r)
BBC Radio 4 FM|1463924700|The Listening Project|||0|0||Omnibus. Fi Glover introduces conversations about art and punctuation, living with MS, and recovering from a stroke.(r)
BBC Radio 4 FM|1463925600|Dangerous Visions: Brave New World|||0|0||Part one of two. Jonathan Holloway's dramatisation of Aldous Huxley's sci-fi novel about a corrupted, hedonistic society where eugenics is practiced as a respected science.
BBC Radio 4 FM|1463929200|Open Book|||0|0||Mariella Frostrup talks to author Kit de Waal about her novel My Name is Leon. Three writers discuss the lengths they went to to ensure factual details in their books were accurate.(r)
BBC Radio 4 FM|1463931000|Poetry Please|||0|0||Roger McGough presents a selection of poetry requests on the theme of wounds and scars, both literal and metaphorical, including works by Hollie McNish, Siegfried Sassoon and Rumi.(r)
BBC Radio 4 FM|1463932800|File on 4|||0|0||Police forces in England and Wales are to get an additional 1,500 firearms officers to help protect the public from terrorism and organised crime. Danny Shaw investigates whether the additional staff will be enough to cope.(r)
BBC Radio 4 FM|1463935200|Profile|||0|0||Friends, adversaries, colleagues and confidants provide an insight into the personality and motivation of Ruth Davidson, leader of the Scottish Conservatives. Mark Coles presents.(r)
BBC Radio 4 FM|1463936040|Shipping Forecast|||0|0||
BBC Radio 4 FM|1463936220|Weather|||0|0||
BBC Radio 4 FM|1463936400|Six O'Clock News|||0|0||
BBC Radio 4 FM|1463937300|Pick of the Week|||0|0||John Waite selects his highlights of the past seven days' radio programmes, including the story of an Irish musical genius and little-known facts about Florence Nightingale.(r)
BBC Radio 4 FM|1463940000|The Archers|||0|0||Rob is having trouble getting through, and Ursula is pleasantly surprised.(r)
BBC Radio 4 FM|1463940900|The Write Stuff|||0|0||James Walton hosts the literary quiz, this week on the English poet William Blake, with captains Sebastian Faulks and John Walsh in attendance alongside guests John O'Farrell and Jane Thynne.(r)
BBC Radio 4 FM|1463942700|Dangerous Visions: Dark Vignettes|||0|0||New series. Short stories presenting disturbing visions of the future. Nicola Walker reads Blackout by Julian Simpson, in which a woman watches order collapse in her city.
BBC Radio 4 FM|1463943600|Feedback|||0|0||Roger Bolton hears listener concerns about the timing of Radio 4's World on the Move day during the EU Referendum. Plus, Soul Music brings back childhood memories and there's discussion about the end of What the Papers Say. ADDRESS: Feedback, PO Box 67234, London SE1P 4AX; phone: 0333 344 4544; e-mail: feedback@bbc.co.uk.(r)
BBC Radio 4 FM|1463945400|Last Word|||0|0||Matthew Bannister pays tribute to animal biomechanics expert Professor Robert McNeill Alexander, Australian TV producer Reg Grundy, and British Elle magazine editor Sally Brampton.(r)
BBC Radio 4 FM|1463947200|Money Box|||0|0||Paul Lewis visits a gold bullion dealer, and considers whether new initiatives go far enough in prompting banks to treat customers better.(r)
BBC Radio 4 FM|1463948760|Radio 4 Appeal|||0|0||Ian McEwan presents an appeal on behalf of SolarAid.(r)
BBC Radio 4 FM|1463949000|In Business|||0|0||Amid concerns about the future of the Port Talbot steelworks and its workers, Peter Day examines the history of the industry in Britain. To find out what went wrong, he hears stories from Port Talbot now and delves into the archive to hear from the heyday of British steel, a time when manufacturing dominated the economy.(r)
BBC Radio 4 FM|1463950740|Weather|||0|0||
BBC Radio 4 FM|1463950800|The Westminster Hour|||0|0||Political magazine, with Carolyn Quinn.(r)
BBC Radio 4 FM|1463954400|The Film Programme|||0|0||Tom Hanks talks about A Hologram for the King and Hollywood's relationship with China, and reveals the advice he was given to have a hit film in the People's Republic.(r)
BBC Radio 4 FM|1463956200|Something Understood|||0|0||Mark Tully examines deterrence, revealing how it often fails to work and can have harmful consequences by preventing people from pursuing other options.(r)
BBC Radio 4 FM|1463958000|News and Weather|||0|0||
BBC Radio 4 FM|1463958900|Thinking Allowed|||0|0||Laurie Taylor examines Glasgow and Russian gangs, including their origins, organisation and meaning in two strikingly different cultures.(r)
BBC Radio 4 FM|1463960700|Bells on Sunday|||0|0||The morning bells from the Parish Church of St Thomas in Hazel Grove, Stockport, ringing Cambridge Surprise Major.(r)
BBC Radio 4 FM|1463960880|Shipping Forecast|||0|0||
BBC Radio 4 FM|1463961600|As BBC World Service|||0|0||
BBC Radio 4 FM|1463977200|Shipping Forecast|||0|0||
BBC Radio 4 FM|1463977800|News Briefing|||0|0||
BBC Radio 4 FM|1463978580|Prayer for the Day|||0|0||Spiritual reflection to start the day with the Very Rev John Chalmers, the former moderator of the Church of Scotland's General Assembly.(r)
BBC Radio 4 FM|1463978700|Farming Today|||0|0||Does the pressure to produce cheap meat fuel the rise in antibiotic resistant superbugs? Tom Heap tells Charlotte Smith about his investigations for tonight's Panorama.(r)
BBC Radio 4 FM|1463979480|Tweet of the Day|||0|0||David Attenborough presents the sound of the pied flycatcher, which travel from Africa to the UK in time for the spring.(r)
BBC Radio 4 FM|1463979600|Today|||0|0||News headlines and sport, presented by Nick Robinson and Sarah Montague. 6.25, 7.25, 8.25 Sports News. 7.48 Thought for the Day with the Rev Dr Jane Leach.(r)
BBC Radio 4 FM|1463990400|Start the Week|||0|0||Andrew Marr is joined by poet Simon Armitage, artist Cornelia Parker, archaeologist Cyprian Broodbank and British Museum curator Aurelia Masson-Berghoff.(r)
BBC Radio 4 FM|1463993100|In the Bonesetter's Waiting Room|||0|0||By Aarathi Prasad, abridged by Pete Nichols. The geneticist and author explores the ancient and modern in Indian medicine, beginning with its seven officials types. Read by Sudha Bhuchar.(r)
BBC Radio 4 FM|1463994000|Woman's Hour|||0|0||Discussion and interviews, presented by Jane Garvey, with Toni Myers. Including at 10.45 the 15 Minute Drama: Part one of Tales of the City: Mary Ann in Autumn, by Armistead Maupin.(r)
BBC Radio 4 FM|1463997600|The Untold|||0|0||Grace Dent follows the story of Mandy Harmon, who was shocked to discover how much the funeral for ex-husband was going to cost and was determined to help her three children with the cost.(r)
BBC Radio 4 FM|1463999400|Fags, Mags and Bags|||0|0||Malcolm and Ramesh's relationship steps up a gear, while Dave dips his toes into the delight of online dating apps. Comedy, written by and starring Sanjeev Kohli and Donald McLeary, with Mina Anwar.(r)
BBC Radio 4 FM|1464001200|News|||0|0||
BBC Radio 4 FM|1464001440|Home Front|||0|0||By Richard Monks. On this day in 1916, the Devon and Exeter Gazette advertised the training of women in the lighter branches of farm work. Meanwhile, Lord Colville takes his daughter to the theatre. Drama set 100 years ago, starring Anton Lesser.(r)
BBC Radio 4 FM|1464002100|You and Yours|||0|0||Consumer and public interest reports.(r)
BBC Radio 4 FM|1464004620|Weather|||0|0||
BBC Radio 4 FM|1464004800|The World at One|||0|0||Analysis of current affairs reports.(r)
BBC Radio 4 FM|1464007500|England: Made in the Middle|||0|0||New series. Helen Castor examines the role of the Anglo-Saxon kingdom of Mercia in the creation of England, asking whether Offa was a greater king than Alfred the Great.
BBC Radio 4 FM|1464008400|The Archers|||0|0||Rob is having trouble getting through, and Ursula is pleasantly surprised.(r)
BBC Radio 4 FM|1464009300|Dangerous Visions|||0|0||By Joseph Wilde. Zenith Genomics seems to offer the ideal solution for a couple unable to have a baby naturally - a perfect, bespoke child. Laura dos Santos and Joseph Kloska star.(r)
BBC Radio 4 FM|1464012000|The 3rd Degree|||0|0||Three undergraduates from the University of Chester challenge their lecturers as Steve Punt hosts another round of the academic quiz show, with specialist subjects including archaeology, English and computer science.(r)
BBC Radio 4 FM|1464013800|The Food Programme|||0|0||The first of two programmes in which author Diana Henry talks to Sheila Dillon about the writers who shaped her passion for food. With readings by Rebecca Ripley and Sam Woolf.(r)
BBC Radio 4 FM|1464015600|Spanish Steps|||0|0||Chris Stewart, author of the best selling Driving Over Lemons, searches for the authentic sound of flamenco, visiting the streets of Granada to uncover its dark past.(r)
BBC Radio 4 FM|1464017400|Beyond Belief|||0|0||Ernie Rea and guests discuss the legacy of the doctrine of original sin.(r)
BBC Radio 4 FM|1464019200|PM|||0|0||Analysis of news headlines, presented by Eddie Mair.(r)
BBC Radio 4 FM|1464022620|Weather|||0|0||
BBC Radio 4 FM|1464022800|Six O'Clock News|||0|0||
BBC Radio 4 FM|1464024480|Referendum Campaign Broadcast|||0|0||By the Vote Leave campaign.(r)
BBC Radio 4 FM|1464024600|Just a Minute|||0|0||Paul Merton, Josie Lawrence, Alexei Sayle and Graham Norton try to speak for 60 seconds without hesitation, repetition or deviation on the panel show chaired by Nicholas Parsons.(r)
BBC Radio 4 FM|1464026400|The Archers|||0|0||Helen cannot relax and Kirsty accepts an apology.(r)
BBC Radio 4 FM|1464027300|Front Row|||0|0||A round-up of arts news and reviews.(r)
BBC Radio 4 FM|1464029100|Tales of the City|||0|0||Lin Coghlan's dramatisation of the eighth instalment of Armistead Maupin's series of novels set in San Francisco. It is 2008 and Mary Anne returns to San Francisco with some big news to share with Michael. Laurel Lefkow stars. Broadcast earlier as part of Woman's Hour.(r)
BBC Radio 4 FM|1464030000|Born in Bradford|||0|0||Winifred Robinson reports on a health study in the West Yorkshire city that has been tracking the fortunes of 14,000 babies from birth over the past seven years.(r)
BBC Radio 4 FM|1464031800|Analysis|||0|0||New series. The return of the programme examining the ideas and forces shaping public policy in Britain and abroad. Linda Pressly asks if being non-binary breaks the last identity taboo, and explores the challenges it creates for the law, society and conventional concepts about gender.(r)
BBC Radio 4 FM|1464033600|The Power of Cute|||0|0||Lucy Cooke explores the biology behind peoples' seeming obsession with all things classed as adorable, and investigates if there is a science to being cute.(r)
BBC Radio 4 FM|1464035400|Start the Week|||0|0||Andrew Marr is joined by poet Simon Armitage, artist Cornelia Parker, archaeologist Cyprian Broodbank and British Museum curator Aurelia Masson-Berghoff.(r)
BBC Radio 4 FM|1464037140|Weather|||0|0||
BBC Radio 4 FM|1464037200|The World Tonight|||0|0||International news round-up.(r)
BBC Radio 4 FM|1464039900|The Bricks That Built the Houses|||0|0||By Kate Tempest. Harry, Becky and Leon flee London with a suitcase full of cash, leaving behind jealous boyfriends, dead-end jobs and irate drug dealers. Read by the author.(r)
BBC Radio 4 FM|1464040800|Don't Make Me Laugh|||0|0||Comedy panel show, hosted by David Baddiel, in which celebrities go against their natural instincts to try not to make an audience laugh. Panellists are Danny Baker, Ross Noble, Mark Watson and Felicity Ward.(r)
BBC Radio 4 FM|1464042600|Today in Parliament|||0|0||Sean Curran presents news, views and analysis of the day's developments in Westminster.(r)
BBC Radio 4 FM|1464044400|News and Weather|||0|0||
BBC Radio 4 FM|1464046200|In the Bonesetter's Waiting Room|||0|0||By Aarathi Prasad, abridged by Pete Nichols. The geneticist and author explores the ancient and modern in Indian medicine, beginning with its seven officials types. Read by Sudha Bhuchar.(n)
BBC Radio 4 FM|1464047280|Shipping Forecast|||0|0||
BBC Radio 4 FM|1464048000|As BBC World Service|||0|0||
BBC Radio 4 FM|1464063600|Shipping Forecast|||0|0||
BBC Radio 4 FM|1464064200|News Briefing|||0|0||
BBC Radio 4 FM|1464064980|Prayer for the Day|||0|0||Spiritual reflection to start the day with the Very Rev John Chalmers, the former moderator of the Church of Scotland's General Assembly.(n)
BBC Radio 4 FM|1464065100|Farming Today|||0|0||Anna Hill presents the latest news about food, farming and the countryside.(n)
BBC Radio 4 FM|1464065880|Tweet of the Day|||0|0||Chris Packham introduces the song of the grey wagtail, a species which tends to nest near flowing water.(n)
BBC Radio 4 FM|1464066000|Today|||0|0||News headlines and sport, presented by John Humphrys and Mishal Husain. 6.25, 7.25, 8.25 Sports News. 6.45 Yesterday in Parliament. 7.48 Thought for the Day, with Anne Atkins.(n)
BBC Radio 4 FM|1464076800|Europeans - The Roots of Identity|||0|0||Historian Margaret MacMillan visits Amsterdam, exploring how a place bound to the sea and the globe developed its idea of Europe. Last in the series.(n)
BBC Radio 4 FM|1464078600|The Ideas That Make Us|||0|0||Bettany Hughes considers the concept of virtue in her study of philosophy, and travels to Athens, Greece, to see how the idea was born and evolved. She meets philosopher Angie Hobbs and the former Greek deputy finance minister Petros Doukas to explore how the notion has been moulded by history, and how modern society has been shaped by it. Last in the series.(n)
BBC Radio 4 FM|1464079500|In the Bonesetter's Waiting Room|||0|0||By Aarathi Prasad, abridged by Pete Nichols. The geneticist explores Indian medicine, continuing with a visit to the shrine of Subawa. Read by Sudha Bhuchar.(n)
BBC Radio 4 FM|1464080400|Woman's Hour|||0|0||Discussion and interviews, presented by Jane Garvey. Including at 10.45 the 15 Minute Drama: Part two of Tales of the City: Mary Ann in Autumn, by Armistead Maupin.(n)
BBC Radio 4 FM|1464084000|Life Under Glass|||0|0||Claire Prentice discovers how a sideshow doctor at Coney Island's amusement fair changed the course of medical history and helped to save premature babies.(n)
BBC Radio 4 FM|1464085800|Punk, the Pistols and the Provinces|||0|0||Mark Hodkinson looks at the impact of punk rock outside of London and, in particular, in Yorkshire, where the Sex Pistols played their first and last gigs outside the capital.(n)
BBC Radio 4 FM|1464087600|News|||0|0||
BBC Radio 4 FM|1464087840|Home Front|||0|0||By Richard Monks. On this day in 1916, the Union Jack was to be flown from every public building for Empire Day, and Dieter feels increasingly isolated.(n)
BBC Radio 4 FM|1464088500|Call You and Yours|||0|0||Consumer affairs, inviting listeners to offer their experiences. PHONE: 0370 010 0444 (Lines open from 10am) email: youandyours@bbc.co.uk.(n)
BBC Radio 4 FM|1464091020|Weather|||0|0||
BBC Radio 4 FM|1464091200|The World at One|||0|0||Analysis of current affairs reports, presented by Martha Kearney.(n)
BBC Radio 4 FM|1464093900|England: Made in the Middle|||0|0||Historian Helen Castor examines the role of the Midlands in the Industrial Revolution, including the story of the Lunar Society - a group of Midland entrepreneurs, enthusiasts and inventors who met up at a location in or near Birmingham once a month, on the Monday nearest the full moon. The Lunar Society counted among its members many of the most innovative thinkers of a particularly innovative age - major figures of the wider Enlightenment whose individual contributions were at least as significant as those of Voltaire in France, Goethe in Germany, and Benjamin Franklin in the United States.(n)
BBC Radio 4 FM|1464094800|The Archers|||0|0||Helen cannot relax and Kirsty accepts an apology.(n)
BBC Radio 4 FM|1464095700|Dangerous Visions: Your Perfect Summer, On Sale Here|||0|0||Ben Tavassoli, Oliver Chris and Claudie Blakley star in Ed Harris's virtual love story, asking what will happen when VR games can deliver real love.(n)
BBC Radio 4 FM|1464098400|The Kitchen Cabinet|||0|0||Jay Rayner hosts the culinary programme from Durham, with panellists Professor Peter Barham, Rachel McCormack and Rob Owen Brown.(n)
BBC Radio 4 FM|1464100200|Shared Experience|||0|0||Fi Glover talks to three men who have chosen to stay at home looking after their young children, while their wives go out to work.(n)
BBC Radio 4 FM|1464102000|Word of Mouth|||0|0||Michael Rosen talks to author Keith Houston about punctuation symbols and how they came to exist, from the first ones up to new inventions like the interrobang. Last in the series.(n)
BBC Radio 4 FM|1464103800|Great Lives|||0|0||Ann Limb, chair of the Scout Association, nominates George Fox, founder of the Quakers. Presented by Matthew Parris.(n)
BBC Radio 4 FM|1464105600|PM|||0|0||Analysis of news headlines, presented by Eddie Mair.(n)
BBC Radio 4 FM|1464109020|Weather|||0|0||
BBC Radio 4 FM|1464109200|Six O'Clock News|||0|0||
BBC Radio 4 FM|1464110880|Referendum Campaign Broadcast|||0|0||By the Stronger in Europe campaign.(n)
BBC Radio 4 FM|1464111000|Isy Suttie's Love Letters|||0|0||Isy Suttie recounts the tale of George and Louise, set against the backdrop of the Matlock Ceilidh over Christmas and New Year 2014. Last in the series.(n)
BBC Radio 4 FM|1464112800|The Archers|||0|0||It's a big day at Home Farm, and Pip has a visitor.(n)
BBC Radio 4 FM|1464113700|Front Row|||0|0||A round-up news and reviews from the arts world.(n)
BBC Radio 4 FM|1464115500|Tales of the City|||0|0||By Armistead Maupin. Dramatised by Lin Coghlan. Mary Anne begins to adapt to life with Michael and Ben, while Jake meets a new man at Pier 39.(n)
BBC Radio 4 FM|1464116400|File on 4|||0|0||The case of Thomas Bourke, a man who has served 22 years in prison for a double murder, but still maintains he did not commit the crime.(n)
BBC Radio 4 FM|1464118800|In Touch|||0|0||News of interest to blind and partially sighted people, presented by Peter White.(n)
BBC Radio 4 FM|1464120000|All in the Mind|||0|0||Claudia Hammond examines pressing issues in the world of psychiatry and mental health.(n)
BBC Radio 4 FM|1464121800|Europeans - The Roots of Identity|||0|0||Historian Margaret MacMillan visits Amsterdam, exploring how a place bound to the sea and the globe developed its idea of Europe. Last in the series.(n)
BBC Radio 4 FM|1464123540|Weather|||0|0||
BBC Radio 4 FM|1464123600|The World Tonight|||0|0||International news round-up, with Ritula Shah.(n)
BBC Radio 4 FM|1464126300|The Bricks That Build the Houses|||0|0||Written and read by Kate Tempest. Becky still dream of dancing, but her reality involves waitressing by day and giving massages in hotels by night.(n)
BBC Radio 4 FM|1464127200|Spotlight Tonight with Nish Kumar|||0|0||The presenter discusses the week's most talked about news items, taking an in-depth look at the biggest stories to scrutinise what is actually going on beneath the bluster.(n)
BBC Radio 4 FM|1464129000|Today in Parliament|||0|0||Susan Hulme presents news, views and analysis of the day's developments in Westminster.(n)
BBC Radio 4 Extra|1463871600|The Turn of the Screw|||0|0||A governess suspects her two charges are harbouring a secret - but the truth may be more terrifying than she could ever have imagined. Neville Teller's dramatisation of Henry James' chilling tale, with Cathy Sara, Joseph Tremain, Lulu Popplewell, Tina Gray and Robert Lister. Originally broadcast in 2004.(r)
BBC Radio 4 Extra|1463875200|Tales of the City|||0|0||Parts 1-5/5. Lin Coghlan's dramatisation of Armistead Maupin's seventh instalment of his series of novels set in San Francisco. It is 2005 and Michael's wedded bliss is interrupted by an unexpected phone call from his brother, while Brian makes plans for the future. Trevor White and Simon Lee Phillips star.(r)
BBC Radio 4 Extra|1463879400|Inheritance Tracks|||0|0||Singer Rick Astley chooses That's Amore, as performed by Dean Martin, and Buck Rogers by Feeder.(r)
BBC Radio 4 Extra|1463879700|Frankly Speaking|||0|0||Room at the Top author John Braine answers the questions in this edition of the BBC Home Service's interview series. First broadcast in 1959.(r)
BBC Radio 4 Extra|1463881500|Could Do Better|||0|0||Robert Booth summons humorist Alan Coren for a quiet word about his school reports. From 1988.(r)
BBC Radio 4 Extra|1463882400|Freud v Jung|||0|0||Lisa Appignanesi delves into the turbulent professional relationship of Sigmund Freud and Carl Jung. She assesses the impact of their work on mankind's understanding of the unconscious mind, and explores how an argument in 1912 drove them apart for good.(r)
BBC Radio 4 Extra|1463886000|The Friend of the Family|||0|0||Chaos erupts in Stepanchikovo, Russia, in 1859, when an ex-sergeant acts as an arbiter of morals and taste. Drama, starring David Suchet. First broadcast December 1984.(r)
BBC Radio 4 Extra|1463891400|Capturing America: Mark Lawson's History of Modern American Literature|||0|0||Writers, including Norman Mailer and Jay McInerney discuss depictions of post-war US foreign policy as America aimed at nipping ideological threats in the bud. They consider EL Doctorow's use of historical parallels, the rise of the espionage thriller, and how the arrival of bloodshed on America's streets with the September 11 attacks changed the mood.
BBC Radio 4 Extra|1463893200|Speaking for Themselves|||0|0||Parts 1-5 of 10. Sylvestra Le Touzel and Alex Jennings read from the personal letters of Clementine and Winston Churchill. Originally broadcast in 1999.(r)
BBC Radio 4 Extra|1463897700|A Woman's World|||0|0||Graham Clarke tells Chris Ledgard about running a WRVS lunch club. The charity - the Women's Royal Voluntary Service - no longer uses its full title and has been taking on male volunteers for many years. Chief executive Lynne Berry discusses the balance between respecting the WRVS's history as a women's organisation, and establishing its new image in the modern world of big charity.(r)
BBC Radio 4 Extra|1463898600|Count Arthur Strong's Radio Show!|||0|0||Comedy drama following the exploits of former variety star Count Arthur Strong. The showbiz veteran tries to reduce his car's insurance premium by proving that Terry Wogan will not be his passenger, causing much confusion along the way. written by and starring Steve Delaney.(r)
BBC Radio 4 Extra|1463900400|Ray's a Laugh|||0|0||Will Ted be able to get over the shock after a new employee arrives? Stars Ted Ray and Kitty Bluett. Originally broadcast in 1958.(r)
BBC Radio 4 Extra|1463902200|Doctor in the House|||0|0||Medic Simon Sparrow's efforts to get a date for the hospital ball turn to chaos. Stars Richard Briers. Originally broadcast in September 1968.(r)
BBC Radio 4 Extra|1463904000|Memories: From Moscow to the Black Sea|||0|0||By Teffi. The Russian writer and satirist's story of how she had to flee her country in the early 1900s. Read by Tracy-Ann Obermann.
BBC Radio 4 Extra|1463908200|Inheritance Tracks|||0|0||Sporty former Spice Girl Melanie C chooses Stevie Wonder's 'I Wish' and 'Eternal Flame' by Bangles.(r)
BBC Radio 4 Extra|1463908500|World Book Club|||0|0||Kate Grenville talks to Harriet Gilbert about her book The Secret River.(r)
BBC Radio 4 Extra|1463912100|The Moth Radio Hour|||0|0||Peter Aguero introduces a special show from New York, with stories about the ties the bind.(r)
BBC Radio 4 Extra|1463914800|Ray's a Laugh|||0|0||Will Ted be able to get over the shock after a new employee arrives? Stars Ted Ray and Kitty Bluett. Originally broadcast in 1958.(r)
BBC Radio 4 Extra|1463916600|Doctor in the House|||0|0||Medic Simon Sparrow's efforts to get a date for the hospital ball turn to chaos. Stars Richard Briers. Originally broadcast in September 1968.(r)
BBC Radio 4 Extra|1463918400|Speaking for Themselves|||0|0||Parts 1-5 of 10. Sylvestra Le Touzel and Alex Jennings read from the personal letters of Clementine and Winston Churchill. Originally broadcast in 1999.(r)
BBC Radio 4 Extra|1463922900|A Woman's World|||0|0||Graham Clarke tells Chris Ledgard about running a WRVS lunch club. The charity - the Women's Royal Voluntary Service - no longer uses its full title and has been taking on male volunteers for many years. Chief executive Lynne Berry discusses the balance between respecting the WRVS's history as a women's organisation, and establishing its new image in the modern world of big charity.(r)
BBC Radio 4 Extra|1463923800|The Typewriter's Tale|||0|0||1907: writer Henry James's typist, Frieda, is drawn to a new arrival at Lamb House in Rye. Read by Sian Thomas.(r)
BBC Radio 4 Extra|1463928300|The Shades of Spring|||0|0||By DH Lawrence. Addy Syson returns to the country of his past in search of the girl he left behind. Peter Meakin reads the short story.(r)
BBC Radio 4 Extra|1463929200|Habakkuk of Ice|||0|0||The story of Second World War inventor Geoffrey Pyke, who designed a battleship made of ice and wood. Fact-based drama by Steve Walker, with Tim McInnerney, Dermot Crowley, Melanie Hudson and Chris Emmett.(r)
BBC Radio 4 Extra|1463932800|Poetry Extra: Paul Celan in Mapesbury Road|||0|0||Writer Toby Litt investigates what compelled master elegist Paul Celan to write a poem about his experience of an ordinary north London street. Along the way, he discovers whom Celan visited while he was there, and asks why such an improbable brief encounter inspired one of the poet's greatest works.
BBC Radio 4 Extra|1463934600|Count Arthur Strong's Radio Show!|||0|0||Comedy drama following the exploits of former variety star Count Arthur Strong. The showbiz veteran tries to reduce his car's insurance premium by proving that Terry Wogan will not be his passenger, causing much confusion along the way. written by and starring Steve Delaney.(r)
BBC Radio 4 Extra|1463936400|Rock of Eye|||0|0||By Anita Sullivan. Three tailors are making a bespoke suit for an up-and-coming politician. The garment has been designed by the mysterious Mrs White, and the fabric they are given seems to change colour and quality along with their moods. As it takes shape, they come to realise the clothing has a powerful effect on anyone who comes into contact with it. Supernatural drama, starring Allan Corduner and Liza Sadovy.(r)
BBC Radio 4 Extra|1463939100|Beware of the Dog|||0|0||On his way back to base following a mission, a badly injured Spitfire pilot is forced to bail out. Read by James Aubrey.(r)
BBC Radio 4 Extra|1463940000|The Moth Radio Hour|||0|0||Peter Aguero introduces a special show from New York, with stories about the ties the bind.(r)
BBC Radio 4 Extra|1463942700|Memories: From Moscow to the Black Sea|||0|0||By Teffi. The Russian writer and satirist's story of how she had to flee her country in the early 1900s. Read by Tracy-Ann Obermann.
BBC Radio 4 Extra|1463946900|Inheritance Tracks|||0|0||Sporty former Spice Girl Melanie C chooses Stevie Wonder's 'I Wish' and 'Eternal Flame' by Bangles.(r)
BBC Radio 4 Extra|1463947200|World Book Club|||0|0||Kate Grenville talks to Harriet Gilbert about her book The Secret River.(r)
BBC Radio 4 Extra|1463950800|Count Arthur Strong's Radio Show!|||0|0||Comedy drama following the exploits of former variety star Count Arthur Strong. The showbiz veteran tries to reduce his car's insurance premium by proving that Terry Wogan will not be his passenger, causing much confusion along the way. written by and starring Steve Delaney.(r)
BBC Radio 4 Extra|1463952600|The Masterson Inheritance|||0|0||Ancient Rome witnesses terror, tyrants and togas. Improvised family saga with Paul Merton and Josie Lawrence. Originally broadcast in June 1994.(r)
BBC Radio 4 Extra|1463954400|John Shuttleworth's Open Mind|||0|0||The Sheffield singer-songwriter tries to solve the Atlantic Ocean mystery. With Sir Robin Knox-Johnston. Originally broadcast in April 2006.(r)
BBC Radio 4 Extra|1463956200|Births, Deaths and Marriages|||0|0||Comedy by and starring David Schneider. Malcolm is distracted by a breast-feeding mother during a birth registration, causing Lorna to believe he may have made his first-ever mistake. With Sarah Hadland and Sandy McDade.(r)
BBC Radio 4 Extra|1463958000|Rock of Eye|||0|0||By Anita Sullivan. Three tailors are making a bespoke suit for an up-and-coming politician. The garment has been designed by the mysterious Mrs White, and the fabric they are given seems to change colour and quality along with their moods. As it takes shape, they come to realise the clothing has a powerful effect on anyone who comes into contact with it. Supernatural drama, starring Allan Corduner and Liza Sadovy.(r)
BBC Radio 4 Extra|1463960700|Beware of the Dog|||0|0||On his way back to base following a mission, a badly injured Spitfire pilot is forced to bail out. Read by James Aubrey.(r)
BBC Radio 4 Extra|1463961600|Speaking for Themselves|||0|0||Parts 1-5 of 10. Sylvestra Le Touzel and Alex Jennings read from the personal letters of Clementine and Winston Churchill. Originally broadcast in 1999.(r)
BBC Radio 4 Extra|1463966100|A Woman's World|||0|0||Graham Clarke tells Chris Ledgard about running a WRVS lunch club. The charity - the Women's Royal Voluntary Service - no longer uses its full title and has been taking on male volunteers for many years. Chief executive Lynne Berry discusses the balance between respecting the WRVS's history as a women's organisation, and establishing its new image in the modern world of big charity.(r)
BBC Radio 4 Extra|1463967000|The Typewriter's Tale|||0|0||1907: writer Henry James's typist, Frieda, is drawn to a new arrival at Lamb House in Rye. Read by Sian Thomas.(r)
BBC Radio 4 Extra|1463971500|The Shades of Spring|||0|0||By DH Lawrence. Addy Syson returns to the country of his past in search of the girl he left behind. Peter Meakin reads the short story.(r)
BBC Radio 4 Extra|1463972400|Habakkuk of Ice|||0|0||The story of Second World War inventor Geoffrey Pyke, who designed a battleship made of ice and wood. Fact-based drama by Steve Walker, with Tim McInnerney, Dermot Crowley, Melanie Hudson and Chris Emmett.(r)
BBC Radio 4 Extra|1463976000|Poetry Extra: Paul Celan in Mapesbury Road|||0|0||Writer Toby Litt investigates what compelled master elegist Paul Celan to write a poem about his experience of an ordinary north London street. Along the way, he discovers whom Celan visited while he was there, and asks why such an improbable brief encounter inspired one of the poet's greatest works.
BBC Radio 4 Extra|1463977800|Count Arthur Strong's Radio Show!|||0|0||Comedy drama following the exploits of former variety star Count Arthur Strong. The showbiz veteran tries to reduce his car's insurance premium by proving that Terry Wogan will not be his passenger, causing much confusion along the way. written by and starring Steve Delaney.(r)
BBC Radio 4 Extra|1463979600|Lord Peter Wimsey - The Nine Tailors|||0|0||The sleuth identifies the body, but he has yet to name the killer. Murder mystery by Dorothy L Sayers, with Ian Carmichael and John Westbrook. Originally broadcast in 1980.(r)
BBC Radio 4 Extra|1463981400|Grayson Perry on Creativity and Imagination|||0|0||Turner Prize-winning ceramicist Grayson Perry sets out to discover what it means to be creative, exposing some of the myths that surround the concept and exploring how the imagination works. Includes contributions by writers Terry Pratchett and Rose Tremain, fashion designer Hussein Chalayan and cultural commentator Stephen Bayley.(r)
BBC Radio 4 Extra|1463983200|Elephants to Catch Eels|||0|0||Tamsyn tries to keep her love-life out of the scandal rags. Comedy, with Lucy Speed, John Bowe, Andrew McGibbon, Cameron Stewart, Martin Hyder and Mark Felgate. First aired in 2003.(r)
BBC Radio 4 Extra|1463985000|Just a Minute|||0|0||The comedy panel show returns for its 75th series, with Paul Merton, John Finnemore, Gyles Brandreth and Sheila Hancock joining host Nicholas Parsons as they try to speak on a given topic for 60 seconds without hesitation, repetition or deviation.(r)
BBC Radio 4 Extra|1463986800|Parsley Sidings|||0|0||Horace decides to restore his grandfather's old train, the Josiah Hepplewhite Rocket, ready for a special exhibition. Comedy, starring Arthur Lowe and Kenneth Connor. First aired in 1972.(r)
BBC Radio 4 Extra|1463988600|J Kingston Platt's Showbiz Handbook|||0|0||The veteran actor recounts a disastrous TV adaptation and its American backer. Comedy, written and performed by Peter Jones. First aired in 1986.(r)
BBC Radio 4 Extra|1463990400|The Write Stuff|||0|0||James Walton hosts the light-hearted literary quiz, with Jane Thynne and Christopher Brookmyre joining captains Lynne Truss and John Walsh. The author is John Donne and the reader Beth Chalmers. First broadcast in 2010.(r)
BBC Radio 4 Extra|1463992200|Tony's|||0|0||The barber's mother threatens to interfere in his unpromising love life. Comedy, with Victor Spinetti, Deborah Watling, John Laurie and Norma Ronald. First aired in 1979.(r)
BBC Radio 4 Extra|1463994000|The Brothers Karamazov|||0|0||In 1880s Russia, the unpredictable Fyodor Karamazov and his sons are re-united to discuss Dmitry's inheritance. Melissa Murray's dramatisation of Fyodor Dostoyevsky's novel, with Roy Marsden, Paul Hilton, Nicholas Boulton, Carl Prekopp and Rachel Atkins. First aired in 2006.(r)
BBC Radio 4 Extra|1463997600|The Human Cradle|||0|0||Saba. By Sulaiman Addonia. The first of three stories by writers from Eritrea, Ethiopia and Somalia on the Horn of Africa. A former cinema employee decides to put on his own screenings inside a refugee camp. Read by Abukar Osman.(r)
BBC Radio 4 Extra|1463998500|Keeping Anne-Marie|||0|0||A woman offers to help her friends by acting as a surrogate mother, but her good intentions backfire when nine months later she changes her mind. Drama by Dave Sheasby, with Geoffrey Whitehead, Hannah Storey, Carolyn Pickles and Sean Baker. Originally broadcast in 2003.(r)
BBC Radio 4 Extra|1464001200|Parsley Sidings|||0|0||Horace decides to restore his grandfather's old train, the Josiah Hepplewhite Rocket, ready for a special exhibition. Comedy, starring Arthur Lowe and Kenneth Connor. First aired in 1972.(r)
BBC Radio 4 Extra|1464003000|J Kingston Platt's Showbiz Handbook|||0|0||The veteran actor recounts a disastrous TV adaptation and its American backer. Comedy, written and performed by Peter Jones. First aired in 1986.(r)
BBC Radio 4 Extra|1464004800|Lord Peter Wimsey - The Nine Tailors|||0|0||The sleuth identifies the body, but he has yet to name the killer. Murder mystery by Dorothy L Sayers, with Ian Carmichael and John Westbrook. Originally broadcast in 1980.(r)
BBC Radio 4 Extra|1464006600|Grayson Perry on Creativity and Imagination|||0|0||Turner Prize-winning ceramicist Grayson Perry sets out to discover what it means to be creative, exposing some of the myths that surround the concept and exploring how the imagination works. Includes contributions by writers Terry Pratchett and Rose Tremain, fashion designer Hussein Chalayan and cultural commentator Stephen Bayley.(r)
BBC Radio 4 Extra|1464008400|The Secret River|||0|0||Ron Cook reads from Kate Grenville's novel about a man transported to Australia in 1806.(r)
BBC Radio 4 Extra|1464009300|In Search of Ourselves: A History of Psychology and the Mind|||0|0||Martin Sixsmith considers how the work of philosopher John Locke and scientist Luigi Galvani, and some of their contemporaries, helped to build the foundations of experimental psychology. The presenter also examines popular fields of study in Victorian times, such as phrenology and physiognomy, and goes behind the scenes at the Science Museum with curator Philip Loring.
BBC Radio 4 Extra|1464010200|Speaking for Themselves|||0|0||Away at war, Churchill writes to Clementine stating he wants to return home early. Sylvestra Le Touzel and Alex Jennings read from the personal letters of Clementine and Winston Churchill. First broadcast in 1999.(r)
BBC Radio 4 Extra|1464011100|How Shall I Tell the Dog?|||0|0||Michael Palin reads from Miles Kington's book written while the columnist was suffering from pancreatic cancer. First aired in 2008.(r)
BBC Radio 4 Extra|1464012000|The Brothers Karamazov|||0|0||In 1880s Russia, the unpredictable Fyodor Karamazov and his sons are re-united to discuss Dmitry's inheritance. Melissa Murray's dramatisation of Fyodor Dostoyevsky's novel, with Roy Marsden, Paul Hilton, Nicholas Boulton, Carl Prekopp and Rachel Atkins. First aired in 2006.(r)
BBC Radio 4 Extra|1464015600|The Write Stuff|||0|0||James Walton hosts the light-hearted literary quiz, with Jane Thynne and Christopher Brookmyre joining captains Lynne Truss and John Walsh. The author is John Donne and the reader Beth Chalmers. First broadcast in 2010.(r)
BBC Radio 4 Extra|1464017400|Tony's|||0|0||The barber's mother threatens to interfere in his unpromising love life. Comedy, with Victor Spinetti, Deborah Watling, John Laurie and Norma Ronald. First aired in 1979.(r)
BBC Radio 4 Extra|1464019200|Elephants to Catch Eels|||0|0||Tamsyn tries to keep her love-life out of the scandal rags. Comedy, with Lucy Speed, John Bowe, Andrew McGibbon, Cameron Stewart, Martin Hyder and Mark Felgate. First aired in 2003.(r)
BBC Radio 4 Extra|1464021000|Just a Minute|||0|0||The comedy panel show returns for its 75th series, with Paul Merton, John Finnemore, Gyles Brandreth and Sheila Hancock joining host Nicholas Parsons as they try to speak on a given topic for 60 seconds without hesitation, repetition or deviation.(r)
BBC Radio 4 Extra|1464022800|The Man Who Was Thursday|||0|0||Gabriel Syme is chased through London's snow to St Paul's by the strange figure of the Professor. Geoffrey Palmer reads from GK Chesterton's chilling tale.(r)
BBC Radio 4 Extra|1464024600|A Good Read|||0|0||Rosie Boycott is joined by Jane Asher and Monty Don to discuss books by Joe Simpson, Adam Nicholson and Christ Stewart. First broadcast in 2002.(r)
BBC Radio 4 Extra|1464026400|Parsley Sidings|||0|0||Horace decides to restore his grandfather's old train, the Josiah Hepplewhite Rocket, ready for a special exhibition. Comedy, starring Arthur Lowe and Kenneth Connor. First aired in 1972.(r)
BBC Radio 4 Extra|1464028200|J Kingston Platt's Showbiz Handbook|||0|0||The veteran actor recounts a disastrous TV adaptation and its American backer. Comedy, written and performed by Peter Jones. First aired in 1986.(r)
BBC Radio 4 Extra|1464030000|Lord Peter Wimsey - The Nine Tailors|||0|0||The sleuth identifies the body, but he has yet to name the killer. Murder mystery by Dorothy L Sayers, with Ian Carmichael and John Westbrook. Originally broadcast in 1980.(r)
BBC Radio 4 Extra|1464031800|Grayson Perry on Creativity and Imagination|||0|0||Turner Prize-winning ceramicist Grayson Perry sets out to discover what it means to be creative, exposing some of the myths that surround the concept and exploring how the imagination works. Includes contributions by writers Terry Pratchett and Rose Tremain, fashion designer Hussein Chalayan and cultural commentator Stephen Bayley.(r)
BBC Radio 4 Extra|1464033600|The Human Cradle|||0|0||Saba. By Sulaiman Addonia. The first of three stories by writers from Eritrea, Ethiopia and Somalia on the Horn of Africa. A former cinema employee decides to put on his own screenings inside a refugee camp. Read by Abukar Osman.(r)
BBC Radio 4 Extra|1464034500|Keeping Anne-Marie|||0|0||A woman offers to help her friends by acting as a surrogate mother, but her good intentions backfire when nine months later she changes her mind. Drama by Dave Sheasby, with Geoffrey Whitehead, Hannah Storey, Carolyn Pickles and Sean Baker. Originally broadcast in 2003.(r)
BBC Radio 4 Extra|1464037200|Just a Minute|||0|0||The comedy panel show returns for its 75th series, with Paul Merton, John Finnemore, Gyles Brandreth and Sheila Hancock joining host Nicholas Parsons as they try to speak on a given topic for 60 seconds without hesitation, repetition or deviation.(r)
BBC Radio 4 Extra|1464039000|Kevin Eldon Will See You Now|||0|0||Sketch show written by Kevin Eldon, with additional material by Jason Hazeley, Joel Morris and Toby Davies. This edition features guests including a silly man, former astronaut Neil Armstrong and a hypnotist. Starring Phil Cornwell, Amelia Bullmore and Julia Davis.(r)
BBC Radio 4 Extra|1464040800|The News Quiz Extra|||0|0||Extended edition of the comedy panel show, featuring out-takes, archive clips and behind-the-scenes material.(r)
BBC Radio 4 Extra|1464043500|Singular Women|||0|0||Celia Imrie plays a shy teacher with an unwanted notoriety. Bittersweet comedies about four very different women. From 1997.(r)
BBC Radio 4 Extra|1464044400|The Man Who Was Thursday|||0|0||Gabriel Syme is chased through London's snow to St Paul's by the strange figure of the Professor. Geoffrey Palmer reads from GK Chesterton's chilling tale.(n)
BBC Radio 4 Extra|1464046200|A Good Read|||0|0||Rosie Boycott is joined by Jane Asher and Monty Don to discuss books by Joe Simpson, Adam Nicholson and Christ Stewart. First broadcast in 2002.(n)
BBC Radio 4 Extra|1464048000|Lord Peter Wimsey - The Nine Tailors|||0|0||The sleuth identifies the body, but he has yet to name the killer. Murder mystery by Dorothy L Sayers, with Ian Carmichael and John Westbrook. Originally broadcast in 1980.(n)
BBC Radio 4 Extra|1464049800|Grayson Perry on Creativity and Imagination|||0|0||Turner Prize-winning ceramicist Grayson Perry sets out to discover what it means to be creative, exposing some of the myths that surround the concept and exploring how the imagination works. Includes contributions by writers Terry Pratchett and Rose Tremain, fashion designer Hussein Chalayan and cultural commentator Stephen Bayley.(n)
BBC Radio 4 Extra|1464051600|The Secret River|||0|0||Ron Cook reads from Kate Grenville's novel about a man transported to Australia in 1806.(n)
BBC Radio 4 Extra|1464052500|In Search of Ourselves: A History of Psychology and the Mind|||0|0||Martin Sixsmith considers how the work of philosopher John Locke and scientist Luigi Galvani, and some of their contemporaries, helped to build the foundations of experimental psychology. The presenter also examines popular fields of study in Victorian times, such as phrenology and physiognomy, and goes behind the scenes at the Science Museum with curator Philip Loring.(n)
BBC Radio 4 Extra|1464053400|Speaking for Themselves|||0|0||Away at war, Churchill writes to Clementine stating he wants to return home early. Sylvestra Le Touzel and Alex Jennings read from the personal letters of Clementine and Winston Churchill. First broadcast in 1999.(n)
BBC Radio 4 Extra|1464054300|How Shall I Tell the Dog?|||0|0||Michael Palin reads from Miles Kington's book written while the columnist was suffering from pancreatic cancer. First aired in 2008.(n)
BBC Radio 4 Extra|1464055200|The Brothers Karamazov|||0|0||In 1880s Russia, the unpredictable Fyodor Karamazov and his sons are re-united to discuss Dmitry's inheritance. Melissa Murray's dramatisation of Fyodor Dostoyevsky's novel, with Roy Marsden, Paul Hilton, Nicholas Boulton, Carl Prekopp and Rachel Atkins. First aired in 2006.(n)
BBC Radio 4 Extra|1464058800|The Write Stuff|||0|0||James Walton hosts the light-hearted literary quiz, with Jane Thynne and Christopher Brookmyre joining captains Lynne Truss and John Walsh. The author is John Donne and the reader Beth Chalmers. First broadcast in 2010.(n)
BBC Radio 4 Extra|1464060600|Tony's|||0|0||The barber's mother threatens to interfere in his unpromising love life. Comedy, with Victor Spinetti, Deborah Watling, John Laurie and Norma Ronald. First aired in 1979.(n)
BBC Radio 4 Extra|1464062400|Elephants to Catch Eels|||0|0||Tamsyn tries to keep her love-life out of the scandal rags. Comedy, with Lucy Speed, John Bowe, Andrew McGibbon, Cameron Stewart, Martin Hyder and Mark Felgate. First aired in 2003.(n)
BBC Radio 4 Extra|1464064200|Just a Minute|||0|0||The comedy panel show returns for its 75th series, with Paul Merton, John Finnemore, Gyles Brandreth and Sheila Hancock joining host Nicholas Parsons as they try to speak on a given topic for 60 seconds without hesitation, repetition or deviation.(n)
BBC Radio 4 Extra|1464066000|Lord Peter Wimsey - The Nine Tailors|||0|0||The upper-class sleuth goes snooping to try and establish who killed Geoffrey Deacon - and how. Murder mystery by Dorothy L Sayers, with Ian Carmichael. Originally broadcast in 1980.(n)
BBC Radio 4 Extra|1464067800|Grayson on His Bike|||0|0||Artist Grayson Perry travels across Bavaria on a highly decorated Kenilworth AM1 motorcycle, accompanied by his teddy bear and childhood hero Alan Measles. Beginning in his home town of Chelmsford, the journey takes Perry via the 1920s Nurburgring racetrack and the Brandhorts Museum of Contemporary Art, before concluding in the town of Backnang, where he delivers a message of goodwill to the local mayor. From 2010.(n)
BBC Radio 4 Extra|1464069600|Linda Smith's A Brief History of Timewasting|||0|0||With London house prices going stratospheric in the East End, Linda gets a valuation. With Jeremy Hardy. First aired in 2002.(n)
BBC Radio 4 Extra|1464071400|Isy Suttie's Love Letters|||0|0||The comedy actress's account of love stories affecting people she has known throughout her life, related through words and song, and accompanied by her guitar. In the third episode, Isy recounts the tale of `The Crank', a Matlock oddball who helped her study the Welsh language. Along the way, Isy picks up a bit of Morse code.(n)
BBC Radio 4 Extra|1464073200|Round the Horne|||0|0||Crofter Kenneth Horne meets Bona Prince Charlie - and bona advertising with Julian and Sandy. With Hugh Paddick. From June 1968.(n)
BBC Radio 4 Extra|1464075000|The Men from the Ministry|||0|0||Confusion, and an ancient Egyptian queen, rule. Stars Deryck Guyler and Richard Murdoch. From July 1974.(n)
BBC Radio 4 Extra|1464076800|The News Quiz Extra|||0|0||Extended edition of the comedy panel show, featuring out-takes, archive clips and behind-the-scenes material.(n)
BBC Radio 4 Extra|1464079500|Singular Women|||0|0||Celia Imrie plays a shy teacher with an unwanted notoriety. Bittersweet comedies about four very different women. From 1997.(n)
BBC Radio 4 Extra|1464080400|The Brothers Karamazov|||0|0||Alyosha attends the bedside of the dying Elder, while the conflict between Dmitry and his father deepens further. Melissa Murray's dramatisation of Fyodor Dostoyevsky's novel, with Roy Marsden, Paul Hilton, Nicholas Boulton, Carl Prekopp and Rachel Atkins. From 2006.(n)
BBC Radio 4 Extra|1464084000|The Human Cradle|||0|0||The Invisible Map, by Maaza Mengiste. An Ethiopian woman who hopes to find a better life in Europe becomes trapped in a Libyan prison. The second of three stories by writers from Eritrea, Ethiopia and Somalia on the Horn of Africa. Read by Adjoa Andoh. From 2012.(n)
BBC Radio 4 Extra|1464084900|Tommies|||0|0||By Nick Warburton. Mickey Bliss returns to the front line as a newly-trained officer, but the Allies are still where they were before the start of the battle of Loos. Drama illustrating the events of a real day at war, exactly 100 years ago to the day, based on eyewitness accounts of the action. From 2015.(n)
BBC Radio 4 Extra|1464087600|Round the Horne|||0|0||Crofter Kenneth Horne meets Bona Prince Charlie - and bona advertising with Julian and Sandy. With Hugh Paddick. From June 1968.(n)
BBC Radio 4 Extra|1464089400|The Men from the Ministry|||0|0||Confusion, and an ancient Egyptian queen, rule. Stars Deryck Guyler and Richard Murdoch. From July 1974.(n)
BBC Radio 4 Extra|1464091200|Lord Peter Wimsey - The Nine Tailors|||0|0||The upper-class sleuth goes snooping to try and establish who killed Geoffrey Deacon - and how. Murder mystery by Dorothy L Sayers, with Ian Carmichael. Originally broadcast in 1980.(n)
BBC Radio 4 Extra|1464093000|Grayson on His Bike|||0|0||Artist Grayson Perry travels across Bavaria on a highly decorated Kenilworth AM1 motorcycle, accompanied by his teddy bear and childhood hero Alan Measles. Beginning in his home town of Chelmsford, the journey takes Perry via the 1920s Nurburgring racetrack and the Brandhorts Museum of Contemporary Art, before concluding in the town of Backnang, where he delivers a message of goodwill to the local mayor. From 2010.(n)
BBC Radio 4 Extra|1464094800|The Secret River|||0|0||Will Thornhill's comfortable life in London with his wife is disturbed when fate intervenes. Ron Cook reads from Kate Grenville's novel. From 2006.(n)
BBC Radio 4 Extra|1464095700|In Search of Ourselves: A History of Psychology and the Mind|||0|0||Martin Sixsmith explores how medical research identified different areas of the brain, and looks at how new ways to measure time aided psychologists assessing the speed of thought. Plus, archivist Subhadra Das explains the impact Francis Galton's statistical mass observations had on psychology. From 2014.(n)
BBC Radio 4 Extra|1464096600|Speaking for Themselves|||0|0||Sylvestra Le Touzel and Alex Jennings read from the personal letters of Clementine and Winston Churchill. From 1999.(n)
BBC Radio 4 Extra|1464097500|How Shall I Tell the Dog?|||0|0||Michael Palin reads from Miles Kington's book written while the columnist was suffering from pancreatic cancer. From 2008.(n)
BBC Radio 4 Extra|1464098400|The Brothers Karamazov|||0|0||Alyosha attends the bedside of the dying Elder, while the conflict between Dmitry and his father deepens further. Melissa Murray's dramatisation of Fyodor Dostoyevsky's novel, with Roy Marsden, Paul Hilton, Nicholas Boulton, Carl Prekopp and Rachel Atkins. From 2006.(n)
BBC Radio 4 Extra|1464102000|Counterpoint|||0|0||Ned Sherrin hosts the music quiz, with Graham Bennett of Surbiton, Jerry Knowles of Selsey and Andrew Taylor from Cambridge. From 2005.(n)
BBC Radio 4 Extra|1464103800|Flying the Flag|||0|0||A diplomatic visit sees the ambassador mix the oil and water of artistic détente. Stars Dinsdale Landen. From December 1990.(n)
BBC Radio 4 Extra|1464105600|Linda Smith's A Brief History of Timewasting|||0|0||With London house prices going stratospheric in the East End, Linda gets a valuation. With Jeremy Hardy. First aired in 2002.(n)
BBC Radio 4 Extra|1464107400|Isy Suttie's Love Letters|||0|0||The comedy actress's account of love stories affecting people she has known throughout her life, related through words and song, and accompanied by her guitar. In the third episode, Isy recounts the tale of `The Crank', a Matlock oddball who helped her study the Welsh language. Along the way, Isy picks up a bit of Morse code.(n)
BBC Radio 4 Extra|1464109200|The Man Who Was Thursday|||0|0||With new-found ally the Professor, Gabriel rests up before they both set off to confront Doctor Bull. Read by Geoffrey Palmer. From 2005.(n)
BBC Radio 4 Extra|1464111000|The Tingle Factor|||0|0||Beatles record producer and composer George Martin talks to Jeremy Nicholas about music which stirs his emotions. From 1992.(n)
BBC Radio 4 Extra|1464112800|Round the Horne|||0|0||Crofter Kenneth Horne meets Bona Prince Charlie - and bona advertising with Julian and Sandy. With Hugh Paddick. From June 1968.(n)
BBC Radio 4 Extra|1464114600|The Men from the Ministry|||0|0||Confusion, and an ancient Egyptian queen, rule. Stars Deryck Guyler and Richard Murdoch. From July 1974.(n)
BBC Radio 4 Extra|1464116400|Lord Peter Wimsey - The Nine Tailors|||0|0||The upper-class sleuth goes snooping to try and establish who killed Geoffrey Deacon - and how. Murder mystery by Dorothy L Sayers, with Ian Carmichael. Originally broadcast in 1980.(n)
BBC Radio 4 Extra|1464118200|Grayson on His Bike|||0|0||Artist Grayson Perry travels across Bavaria on a highly decorated Kenilworth AM1 motorcycle, accompanied by his teddy bear and childhood hero Alan Measles. Beginning in his home town of Chelmsford, the journey takes Perry via the 1920s Nurburgring racetrack and the Brandhorts Museum of Contemporary Art, before concluding in the town of Backnang, where he delivers a message of goodwill to the local mayor. From 2010.(n)
BBC Radio 4 Extra|1464120000|The Human Cradle|||0|0||The Invisible Map, by Maaza Mengiste. An Ethiopian woman who hopes to find a better life in Europe becomes trapped in a Libyan prison. The second of three stories by writers from Eritrea, Ethiopia and Somalia on the Horn of Africa. Read by Adjoa Andoh. From 2012.(n)
BBC Radio 4 Extra|1464120900|Tommies|||0|0||By Nick Warburton. Mickey Bliss returns to the front line as a newly-trained officer, but the Allies are still where they were before the start of the battle of Loos. Drama illustrating the events of a real day at war, exactly 100 years ago to the day, based on eyewitness accounts of the action. From 2015.(n)
BBC Radio 4 Extra|1464123600|Isy Suttie's Love Letters|||0|0||The comedy actress's account of love stories affecting people she has known throughout her life, related through words and song, and accompanied by her guitar. In the third episode, Isy recounts the tale of `The Crank', a Matlock oddball who helped her study the Welsh language. Along the way, Isy picks up a bit of Morse code.(n)
BBC Radio 4 Extra|1464125400|The Guns of Adam Riches|||0|0||The 2011 Edinburgh Award-winning comedian draws inspiration from the Wild West to tell the story of cowboy Big Rich. Comedy offering a selection of fast-paced, offbeat sketches, songs, and audience interaction, with Cariad Lloyd and Jim Johnson. From 2013.(n)
BBC Radio 4 Extra|1464126900|The Comedy Club Interview|||0|0||A chat with a guest from the world of comedy.(n)
BBC Radio 4 Extra|1464127200|Vent|||0|0||Despite his coma, Ben finds the strength to punch his physiotherapist, which Mary and Mum take as a sign of progress. Meanwhile, a winged angel and Elvis Presley haunt the patient's dreams. Comedy, with Neil Pearson, Josie Lawrence, Leslie Ash, Fiona Allen and Dave Lamb. First aired in 2006.(n)
BBC Radio 4 Extra|1464129000|The Wilson Dixon Line|||0|0||Country singer Wilson Dixon recounts how ageing hermit Uncle Wilbour helped him get his life back together after his wife Maureen left him. Humorous songs and anecdotes, written and performed by Jesse Griffin, with Jesse Budd. Originally broadcast in 2009.(n)
BBC Radio 4 LW|1463871600|News and Weather|||0|0||
BBC Radio 4 LW|1463873400|Stories from Songwriters|||0|0||The first in a series of specially commissioned stories by songwriters, beginning with Sunset to Break Your Heart by Barb Jungr - a touching story that is set on the Shetland Islands. Read by Suranne Jones.(r)
BBC Radio 4 LW|1463874480|Shipping Forecast|||0|0||
BBC Radio 4 LW|1463875200|As BBC World Service|||0|0||
BBC Radio 4 LW|1463890800|Shipping Forecast|||0|0||
BBC Radio 4 LW|1463891400|News Briefing|||0|0||
BBC Radio 4 LW|1463892180|Bells on Sunday|||0|0||The morning bells from the Parish Church of St Thomas in Hazel Grove, Stockport, ringing Cambridge Surprise Major.(r)
BBC Radio 4 LW|1463892300|Profile|||0|0||Friends, adversaries, colleagues and confidants provide an insight into the personality and motivation of Ruth Davidson, leader of the Scottish Conservatives. Mark Coles presents.(r)
BBC Radio 4 LW|1463893200|News Headlines|||0|0||
BBC Radio 4 LW|1463893500|Something Understood|||0|0||Mark Tully examines deterrence, revealing how it often fails to work and can have harmful consequences by preventing people from pursuing other options.(r)
BBC Radio 4 LW|1463895300|Living World|||0|0||Archive programme in which Lionel Kelleway tracks down radio-tagged hedgehogs as they wake up from hibernation and enter into courtship rituals. Introduced by Chris Packham.(r)
BBC Radio 4 LW|1463896620|Weather|||0|0||
BBC Radio 4 LW|1463896800|News|||0|0||
BBC Radio 4 LW|1463897220|Sunday Papers|||0|0||Review of the latest news stories making the headlines.(r)
BBC Radio 4 LW|1463897400|Sunday|||0|0||Thomas Becket's relic; a new book giving voice to Transgender Christians and the World Humanitarian Summit, some of the stories in this week's programme.(r)
BBC Radio 4 LW|1463900100|Radio 4 Appeal|||0|0||Ian McEwan presents an appeal on behalf of SolarAid.(r)
BBC Radio 4 LW|1463900220|Weather|||0|0||
BBC Radio 4 LW|1463900400|News|||0|0||
BBC Radio 4 LW|1463900820|Sunday Papers|||0|0||Review of the latest news stories making the headlines.(r)
BBC Radio 4 LW|1463901000|Sunday Worship|||0|0||A Mass for Trinity Sunday live from St Anne's Cathedral, Leeds.(r)
BBC Radio 4 LW|1463903280|A Point of View|||0|0||Will Self questions whether the mind is stronger than the body, and what effect the ubiquity of psychiatrists and psychoanalysts plays in modern Britain.(r)
BBC Radio 4 LW|1463903880|Tweet of the Day|||0|0||Miranda Krestovnikoff presents the unusual chirring sound of the nightjar, a bird often heard calling on summer evenings.(r)
BBC Radio 4 LW|1463904000|Broadcasting House|||0|0||A discussion on the week's major headlines, presented by Paddy O'Connell.(r)
BBC Radio 4 LW|1463907600|The Archers|||0|0||Omnibus. Peggy makes a decision, and there is an awkward moment at the Bull.(c)
BBC Radio 4 LW|1463912100|Desert Island Discs|||0|0||Motown producer Berry Gordy talks to Kirsty Young and selects eight records to take to the mythical island.(c)
BBC Radio 4 LW|1463914800|News Headlines|||0|0||
BBC Radio 4 LW|1463914860|Shipping Forecast|||0|0||
BBC Radio 4 LW|1463915040|Just a Minute|||0|0||The comedy panel show returns for its 75th series, with Paul Merton, John Finnemore, Gyles Brandreth and Sheila Hancock joining host Nicholas Parsons as they try to speak on a given topic for 60 seconds without hesitation, repetition or deviation.(c)
BBC Radio 4 LW|1463916600|The Food Programme|||0|0||The first of two programmes in which author Diana Henry talks to Sheila Dillon about the writers who shaped her passion for food. With readings by Rebecca Ripley and Sam Woolf.(c)
BBC Radio 4 LW|1463918220|Weather|||0|0||
BBC Radio 4 LW|1463918400|The World This Weekend|||0|0||Global news and analysis, presented by Mark Mardell.(c)
BBC Radio 4 LW|1463920200|Jutland: The Battle that Won the War|||0|0||Lord Alan West explains why he believes Jutland was the most important First World War battle, a strategic victory that directly paved the way for allied victory.(c)
BBC Radio 4 LW|1463922000|Gardeners' Question Time|||0|0||Eric Robson hosts a correspondence edition from Ness Botanic Gardens in The Wirral, where Christine Walkden, Bob Flowerdew and Pippa Greenwood answer listeners' queries.(c)
BBC Radio 4 LW|1463924700|The Listening Project|||0|0||Omnibus. Fi Glover introduces conversations about art and punctuation, living with MS, and recovering from a stroke.(c)
BBC Radio 4 LW|1463925600|Dangerous Visions: Brave New World|||0|0||Part one of two. Jonathan Holloway's dramatisation of Aldous Huxley's sci-fi novel about a corrupted, hedonistic society where eugenics is practiced as a respected science.(c)
BBC Radio 4 LW|1463929200|Open Book|||0|0||Mariella Frostrup talks to author Kit de Waal about her novel My Name is Leon. Three writers discuss the lengths they went to to ensure factual details in their books were accurate.(c)
BBC Radio 4 LW|1463931000|Poetry Please|||0|0||Roger McGough presents a selection of poetry requests on the theme of wounds and scars, both literal and metaphorical, including works by Hollie McNish, Siegfried Sassoon and Rumi.(c)
BBC Radio 4 LW|1463932800|File on 4|||0|0||Police forces in England and Wales are to get an additional 1,500 firearms officers to help protect the public from terrorism and organised crime. Danny Shaw investigates whether the additional staff will be enough to cope.(c)
BBC Radio 4 LW|1463935200|Profile|||0|0||Friends, adversaries, colleagues and confidants provide an insight into the personality and motivation of Ruth Davidson, leader of the Scottish Conservatives. Mark Coles presents.(c)
BBC Radio 4 LW|1463936040|Shipping Forecast|||0|0||
BBC Radio 4 LW|1463936220|Weather|||0|0||
BBC Radio 4 LW|1463936400|Six O'Clock News|||0|0||
BBC Radio 4 LW|1463937300|Pick of the Week|||0|0||John Waite selects his highlights of the past seven days' radio programmes, including the story of an Irish musical genius and little-known facts about Florence Nightingale.(c)
BBC Radio 4 LW|1463940000|The Archers|||0|0||Rob is having trouble getting through, and Ursula is pleasantly surprised.(r)
BBC Radio 4 LW|1463940900|The Write Stuff|||0|0||James Walton hosts the literary quiz, this week on the English poet William Blake, with captains Sebastian Faulks and John Walsh in attendance alongside guests John O'Farrell and Jane Thynne.(r)
BBC Radio 4 LW|1463942700|Dangerous Visions: Dark Vignettes|||0|0||New series. Short stories presenting disturbing visions of the future. Nicola Walker reads Blackout by Julian Simpson, in which a woman watches order collapse in her city.
BBC Radio 4 LW|1463943600|Feedback|||0|0||Roger Bolton hears listener concerns about the timing of Radio 4's World on the Move day during the EU Referendum. Plus, Soul Music brings back childhood memories and there's discussion about the end of What the Papers Say. ADDRESS: Feedback, PO Box 67234, London SE1P 4AX; phone: 0333 344 4544; e-mail: feedback@bbc.co.uk.(r)
BBC Radio 4 LW|1463945400|Last Word|||0|0||Matthew Bannister pays tribute to animal biomechanics expert Professor Robert McNeill Alexander, Australian TV producer Reg Grundy, and British Elle magazine editor Sally Brampton.(r)
BBC Radio 4 LW|1463947200|Money Box|||0|0||Paul Lewis visits a gold bullion dealer, and considers whether new initiatives go far enough in prompting banks to treat customers better.(r)
BBC Radio 4 LW|1463948760|Radio 4 Appeal|||0|0||Ian McEwan presents an appeal on behalf of SolarAid.(r)
BBC Radio 4 LW|1463949000|In Business|||0|0||Amid concerns about the future of the Port Talbot steelworks and its workers, Peter Day examines the history of the industry in Britain. To find out what went wrong, he hears stories from Port Talbot now and delves into the archive to hear from the heyday of British steel, a time when manufacturing dominated the economy.(r)
BBC Radio 4 LW|1463950740|Weather|||0|0||
BBC Radio 4 LW|1463950800|The Westminster Hour|||0|0||Political magazine, with Carolyn Quinn.(r)
BBC Radio 4 LW|1463954400|The Film Programme|||0|0||Tom Hanks talks about A Hologram for the King and Hollywood's relationship with China, and reveals the advice he was given to have a hit film in the People's Republic.(r)
BBC Radio 4 LW|1463956200|Something Understood|||0|0||Mark Tully examines deterrence, revealing how it often fails to work and can have harmful consequences by preventing people from pursuing other options.(r)
BBC Radio 4 LW|1463958000|News and Weather|||0|0||
BBC Radio 4 LW|1463958900|Thinking Allowed|||0|0||Laurie Taylor examines Glasgow and Russian gangs, including their origins, organisation and meaning in two strikingly different cultures.(r)
BBC Radio 4 LW|1463960700|Bells on Sunday|||0|0||The morning bells from the Parish Church of St Thomas in Hazel Grove, Stockport, ringing Cambridge Surprise Major.(r)
BBC Radio 4 LW|1463960880|Shipping Forecast|||0|0||
BBC Radio 4 LW|1463961600|As BBC World Service|||0|0||
BBC Radio 4 LW|1463977200|Shipping Forecast|||0|0||
BBC Radio 4 LW|1463977800|News Briefing|||0|0||
BBC Radio 4 LW|1463978580|Prayer for the Day|||0|0||Spiritual reflection to start the day with the Very Rev John Chalmers, the former moderator of the Church of Scotland's General Assembly.(r)
BBC Radio 4 LW|1463978700|Farming Today|||0|0||Does the pressure to produce cheap meat fuel the rise in antibiotic resistant superbugs? Tom Heap tells Charlotte Smith about his investigations for tonight's Panorama.(r)
BBC Radio 4 LW|1463979480|Tweet of the Day|||0|0||David Attenborough presents the sound of the pied flycatcher, which travel from Africa to the UK in time for the spring.(r)
BBC Radio 4 LW|1463979600|Today|||0|0||News headlines and sport, presented by Nick Robinson and Sarah Montague. 6.25, 7.25, 8.25 Sports News. 7.48 Thought for the Day with the Rev Dr Jane Leach.(r)
BBC Radio 4 LW|1463990400|Start the Week|||0|0||Andrew Marr is joined by poet Simon Armitage, artist Cornelia Parker, archaeologist Cyprian Broodbank and British Museum curator Aurelia Masson-Berghoff.(r)
BBC Radio 4 LW|1463993100|Daily Service|||0|0||An act of worship, featuring readings from scripture and a range of choral music, led by the Rev Roger Hutchings. Praise We Now the Word of Grace (Savannah). Galatians 1: 6-12. Let All the World (Dyson). God Has Spoken by His Prophets (Blaenwaern). With Manchester Chamber Choir. Director of Music: Jonathan Lo. Organist: Shaun Turnbull.(r)
BBC Radio 4 LW|1463994000|Woman's Hour|||0|0||Discussion and interviews, presented by Jane Garvey, with Toni Myers. Including at 10.45 the 15 Minute Drama: Part one of Tales of the City: Mary Ann in Autumn, by Armistead Maupin.(c)
BBC Radio 4 LW|1463997600|The Untold|||0|0||Grace Dent follows the story of Mandy Harmon, who was shocked to discover how much the funeral for ex-husband was going to cost and was determined to help her three children with the cost.(c)
BBC Radio 4 LW|1463999400|Fags, Mags and Bags|||0|0||Malcolm and Ramesh's relationship steps up a gear, while Dave dips his toes into the delight of online dating apps. Comedy, written by and starring Sanjeev Kohli and Donald McLeary, with Mina Anwar.(c)
BBC Radio 4 LW|1464001200|News|||0|0||
BBC Radio 4 LW|1464001260|Shipping Forecast|||0|0||
BBC Radio 4 LW|1464001440|Home Front|||0|0||By Richard Monks. On this day in 1916, the Devon and Exeter Gazette advertised the training of women in the lighter branches of farm work. Meanwhile, Lord Colville takes his daughter to the theatre. Drama set 100 years ago, starring Anton Lesser.(c)
BBC Radio 4 LW|1464002100|You and Yours|||0|0||Consumer and public interest reports.(c)
BBC Radio 4 LW|1464004620|Weather|||0|0||
BBC Radio 4 LW|1464004800|The World at One|||0|0||Analysis of current affairs reports.(c)
BBC Radio 4 LW|1464007500|England: Made in the Middle|||0|0||Helen Castor examines the role of the Anglo-Saxon kingdom of Mercia in the creation of England, asking whether Offa was a greater king than Alfred the Great.(c)
BBC Radio 4 LW|1464008400|The Archers|||0|0||Rob is having trouble getting through, and Ursula is pleasantly surprised.(c)
BBC Radio 4 LW|1464009300|Dangerous Visions|||0|0||By Joseph Wilde. Zenith Genomics seems to offer the ideal solution for a couple unable to have a baby naturally - a perfect, bespoke child. Laura dos Santos and Joseph Kloska star.(c)
BBC Radio 4 LW|1464012000|The 3rd Degree|||0|0||Three undergraduates from the University of Chester challenge their lecturers as Steve Punt hosts another round of the academic quiz show, with specialist subjects including archaeology, English and computer science.(c)
BBC Radio 4 LW|1464013800|The Food Programme|||0|0||The first of two programmes in which author Diana Henry talks to Sheila Dillon about the writers who shaped her passion for food. With readings by Rebecca Ripley and Sam Woolf.(c)
BBC Radio 4 LW|1464015600|Spanish Steps|||0|0||Chris Stewart, author of the best selling Driving Over Lemons, searches for the authentic sound of flamenco, visiting the streets of Granada to uncover its dark past.(c)
BBC Radio 4 LW|1464017400|Beyond Belief|||0|0||Ernie Rea and guests discuss the legacy of the doctrine of original sin.(c)
BBC Radio 4 LW|1464019200|PM|||0|0||Analysis of news headlines, presented by Eddie Mair.(c)
BBC Radio 4 LW|1464022440|Shipping Forecast|||0|0||
BBC Radio 4 LW|1464022620|Weather|||0|0||
BBC Radio 4 LW|1464022800|Six O'Clock News|||0|0||
BBC Radio 4 LW|1464024480|Referendum Campaign Broadcast|||0|0||By the Vote Leave campaign.(c)
BBC Radio 4 LW|1464024600|Just a Minute|||0|0||Paul Merton, Josie Lawrence, Alexei Sayle and Graham Norton try to speak for 60 seconds without hesitation, repetition or deviation on the panel show chaired by Nicholas Parsons.(c)
BBC Radio 4 LW|1464026400|The Archers|||0|0||Helen cannot relax and Kirsty accepts an apology.(r)
BBC Radio 4 LW|1464027300|Front Row|||0|0||A round-up of arts news and reviews.(r)
BBC Radio 4 LW|1464029100|Tales of the City|||0|0||Lin Coghlan's dramatisation of the eighth instalment of Armistead Maupin's series of novels set in San Francisco. It is 2008 and Mary Anne returns to San Francisco with some big news to share with Michael. Laurel Lefkow stars. Broadcast earlier as part of Woman's Hour.(r)
BBC Radio 4 LW|1464030000|Born in Bradford|||0|0||Winifred Robinson reports on a health study in the West Yorkshire city that has been tracking the fortunes of 14,000 babies from birth over the past seven years.(r)
BBC Radio 4 LW|1464031800|Analysis|||0|0||New series. The return of the programme examining the ideas and forces shaping public policy in Britain and abroad. Linda Pressly asks if being non-binary breaks the last identity taboo, and explores the challenges it creates for the law, society and conventional concepts about gender.(r)
BBC Radio 4 LW|1464033600|The Power of Cute|||0|0||Lucy Cooke explores the biology behind peoples' seeming obsession with all things classed as adorable, and investigates if there is a science to being cute.(r)
BBC Radio 4 LW|1464035400|Start the Week|||0|0||Andrew Marr is joined by poet Simon Armitage, artist Cornelia Parker, archaeologist Cyprian Broodbank and British Museum curator Aurelia Masson-Berghoff.(r)
BBC Radio 4 LW|1464037140|Weather|||0|0||
BBC Radio 4 LW|1464037200|The World Tonight|||0|0||International news round-up.(r)
BBC Radio 4 LW|1464039900|The Bricks That Built the Houses|||0|0||By Kate Tempest. Harry, Becky and Leon flee London with a suitcase full of cash, leaving behind jealous boyfriends, dead-end jobs and irate drug dealers. Read by the author.(r)
BBC Radio 4 LW|1464040800|Don't Make Me Laugh|||0|0||Comedy panel show, hosted by David Baddiel, in which celebrities go against their natural instincts to try not to make an audience laugh. Panellists are Danny Baker, Ross Noble, Mark Watson and Felicity Ward.(r)
BBC Radio 4 LW|1464042600|Today in Parliament|||0|0||Sean Curran presents news, views and analysis of the day's developments in Westminster.(r)
BBC Radio 4 LW|1464044400|News and Weather|||0|0||
BBC Radio 4 LW|1464046200|In the Bonesetter's Waiting Room|||0|0||By Aarathi Prasad, abridged by Pete Nichols. The geneticist and author explores the ancient and modern in Indian medicine, beginning with its seven officials types. Read by Sudha Bhuchar.(n)
BBC Radio 4 LW|1464047280|Shipping Forecast|||0|0||
BBC Radio 4 LW|1464048000|As BBC World Service|||0|0||
BBC Radio 4 LW|1464063600|Shipping Forecast|||0|0||
BBC Radio 4 LW|1464064200|News Briefing|||0|0||
BBC Radio 4 LW|1464064980|Prayer for the Day|||0|0||Spiritual reflection to start the day with the Very Rev John Chalmers, the former moderator of the Church of Scotland's General Assembly.(n)
BBC Radio 4 LW|1464065100|Farming Today|||0|0||Anna Hill presents the latest news about food, farming and the countryside.(n)
BBC Radio 4 LW|1464065880|Tweet of the Day|||0|0||Chris Packham introduces the song of the grey wagtail, a species which tends to nest near flowing water.(n)
BBC Radio 4 LW|1464066000|Today|||0|0||News headlines and sport, presented by John Humphrys and Mishal Husain. 6.25, 7.25, 8.25 Sports News. 6.45 Yesterday in Parliament. 7.48 Thought for the Day, with Anne Atkins.(n)
BBC Radio 4 LW|1464075060|Yesterday in Parliament|||0|0||Susan Hulme presents an update on the latest political proceedings.(n)
BBC Radio 4 LW|1464076800|Europeans - The Roots of Identity|||0|0||Historian Margaret MacMillan visits Amsterdam, exploring how a place bound to the sea and the globe developed its idea of Europe. Last in the series.(n)
BBC Radio 4 LW|1464078600|The Ideas That Make Us|||0|0||Bettany Hughes considers the concept of virtue in her study of philosophy, and travels to Athens, Greece, to see how the idea was born and evolved. She meets philosopher Angie Hobbs and the former Greek deputy finance minister Petros Doukas to explore how the notion has been moulded by history, and how modern society has been shaped by it. Last in the series.(n)
BBC Radio 4 LW|1464079500|Daily Service|||0|0||Led by John Forrest. Lead Us Heavenly Father, Lead Us. 1 Corinthians 3, vv1-9. When a Knight Won His Spurs (Clarke/Walker), There Is a Higher Throne (Getty).(n)
BBC Radio 4 LW|1464080400|Woman's Hour|||0|0||Discussion and interviews, presented by Jane Garvey. Including at 10.45 the 15 Minute Drama: Part two of Tales of the City: Mary Ann in Autumn, by Armistead Maupin.(n)
BBC Radio 4 LW|1464084000|Life Under Glass|||0|0||Claire Prentice discovers how a sideshow doctor at Coney Island's amusement fair changed the course of medical history and helped to save premature babies.(n)
BBC Radio 4 LW|1464085800|Punk, the Pistols and the Provinces|||0|0||Mark Hodkinson looks at the impact of punk rock outside of London and, in particular, in Yorkshire, where the Sex Pistols played their first and last gigs outside the capital.(n)
BBC Radio 4 LW|1464087600|News|||0|0||
BBC Radio 4 LW|1464087660|Shipping Forecast|||0|0||
BBC Radio 4 LW|1464087840|Home Front|||0|0||By Richard Monks. On this day in 1916, the Union Jack was to be flown from every public building for Empire Day, and Dieter feels increasingly isolated.(n)
BBC Radio 4 LW|1464088500|Call You and Yours|||0|0||Consumer affairs, inviting listeners to offer their experiences. PHONE: 0370 010 0444 (Lines open from 10am) email: youandyours@bbc.co.uk.(n)
BBC Radio 4 LW|1464091020|Weather|||0|0||
BBC Radio 4 LW|1464091200|The World at One|||0|0||Analysis of current affairs reports, presented by Martha Kearney.(n)
BBC Radio 4 LW|1464093900|England: Made in the Middle|||0|0||Historian Helen Castor examines the role of the Midlands in the Industrial Revolution, including the story of the Lunar Society - a group of Midland entrepreneurs, enthusiasts and inventors who met up at a location in or near Birmingham once a month, on the Monday nearest the full moon. The Lunar Society counted among its members many of the most innovative thinkers of a particularly innovative age - major figures of the wider Enlightenment whose individual contributions were at least as significant as those of Voltaire in France, Goethe in Germany, and Benjamin Franklin in the United States.(n)
BBC Radio 4 LW|1464094800|The Archers|||0|0||Helen cannot relax and Kirsty accepts an apology.(n)
BBC Radio 4 LW|1464095700|Dangerous Visions: Your Perfect Summer, On Sale Here|||0|0||Ben Tavassoli, Oliver Chris and Claudie Blakley star in Ed Harris's virtual love story, asking what will happen when VR games can deliver real love.(n)
BBC Radio 4 LW|1464098400|The Kitchen Cabinet|||0|0||Jay Rayner hosts the culinary programme from Durham, with panellists Professor Peter Barham, Rachel McCormack and Rob Owen Brown.(n)
BBC Radio 4 LW|1464100200|Shared Experience|||0|0||Fi Glover talks to three men who have chosen to stay at home looking after their young children, while their wives go out to work.(n)
BBC Radio 4 LW|1464102000|Word of Mouth|||0|0||Michael Rosen talks to author Keith Houston about punctuation symbols and how they came to exist, from the first ones up to new inventions like the interrobang. Last in the series.(n)
BBC Radio 4 LW|1464103800|Great Lives|||0|0||Ann Limb, chair of the Scout Association, nominates George Fox, founder of the Quakers. Presented by Matthew Parris.(n)
BBC Radio 4 LW|1464105600|PM|||0|0||Analysis of news headlines, presented by Eddie Mair.(n)
BBC Radio 4 LW|1464108840|Shipping Forecast|||0|0||
BBC Radio 4 LW|1464109020|Weather|||0|0||
BBC Radio 4 LW|1464109200|Six O'Clock News|||0|0||
BBC Radio 4 LW|1464110880|Referendum Campaign Broadcast|||0|0||By the Stronger in Europe campaign.(n)
BBC Radio 4 LW|1464111000|Isy Suttie's Love Letters|||0|0||Isy Suttie recounts the tale of George and Louise, set against the backdrop of the Matlock Ceilidh over Christmas and New Year 2014. Last in the series.(n)
BBC Radio 4 LW|1464112800|The Archers|||0|0||It's a big day at Home Farm, and Pip has a visitor.(n)
BBC Radio 4 LW|1464113700|Front Row|||0|0||A round-up news and reviews from the arts world.(n)
BBC Radio 4 LW|1464115500|Tales of the City|||0|0||By Armistead Maupin. Dramatised by Lin Coghlan. Mary Anne begins to adapt to life with Michael and Ben, while Jake meets a new man at Pier 39.(n)
BBC Radio 4 LW|1464116400|File on 4|||0|0||The case of Thomas Bourke, a man who has served 22 years in prison for a double murder, but still maintains he did not commit the crime.(n)
BBC Radio 4 LW|1464118800|In Touch|||0|0||News of interest to blind and partially sighted people, presented by Peter White.(n)
BBC Radio 4 LW|1464120000|All in the Mind|||0|0||Claudia Hammond examines pressing issues in the world of psychiatry and mental health.(n)
BBC Radio 4 LW|1464121800|Europeans - The Roots of Identity|||0|0||Historian Margaret MacMillan visits Amsterdam, exploring how a place bound to the sea and the globe developed its idea of Europe. Last in the series.(n)
BBC Radio 4 LW|1464123540|Weather|||0|0||
BBC Radio 4 LW|1464123600|The World Tonight|||0|0||International news round-up, with Ritula Shah.(n)
BBC Radio 4 LW|1464126300|The Bricks That Build the Houses|||0|0||Written and read by Kate Tempest. Becky still dream of dancing, but her reality involves waitressing by day and giving massages in hotels by night.(n)
BBC Radio 4 LW|1464127200|Spotlight Tonight with Nish Kumar|||0|0||The presenter discusses the week's most talked about news items, taking an in-depth look at the biggest stories to scrutinise what is actually going on beneath the bluster.(n)
BBC Radio 4 LW|1464129000|Today in Parliament|||0|0||Susan Hulme presents news, views and analysis of the day's developments in Westminster.(n)
BBC Radio 5 live|1463871600|5 Live in Short|||0|0||Highlights from the past seven days, including the biggest news and sports stories of the week.(r)
BBC Radio 5 live|1463875200|Up All Night|||0|0||With Dotun Adebayo. Including the New York hour, nominations for the Virtual Jukebox and updates from BBC correspondents in cities around the world.(r)
BBC Radio 5 live|1463889600|The Non League Football Show|||0|0||Caroline Barker examines what is good about non-league football from the perspective of the fans.(r)
BBC Radio 5 live|1463893200|Sunday Breakfast|||0|0||Chris Warburton and Sam Walker present the day's main news stories, the latest sport, travel and weather.(r)
BBC Radio 5 live|1463904000|SportsWeek|||0|0||Garry Richardson and guests discuss the past seven days' events.(r)
BBC Radio 5 live|1463907600|Pienaar's Politics|||0|0||John Pienaar shares political observations, with news and interviews from Westminster.(r)
BBC Radio 5 live|1463911200|All About Property with Gabby Logan|||0|0||The sports presenter turns her attention to property, fronting the UK's first radio programme totally dedicated to the subject. She is joined by experts to talk about buying, selling, renting or finding the perfect holiday home.(r)
BBC Radio 5 live|1463914800|5 Live Sport|||0|0||Jonathan Overend introduces football coverage of the Scottish Premiership play-off final second-leg match, French Open tennis and updates of England v Sri Lanka from Headingley.(r)
BBC Radio 5 live|1463931000|5 Live Sport|||0|0||Kelly Cates presents build-up to this afternoon's friendly between England and Turkey.(r)
BBC Radio 5 live|1463933700|5 Live Sport: International Football 2015-16|||0|0||England v Turkey (Kick-off 5.15pm). Commentary on the international friendly at Etihad Stadium in Manchester.
BBC Radio 5 live|1463941800|The 5 Live Hit List|||0|0||Emma Barnett presents a rundown of the top 40 news, politics, sport and showbiz stories of the week, which are making the biggest impact online.(r)
BBC Radio 5 live|1463950800|Stephen Nolan|||0|0||
BBC Radio 5 live|1463961600|Up All Night|||0|0||Dotun Adebayo with the top stories from around the world, including a look at the US papers and the Monday morning phone-in.(r)
BBC Radio 5 live|1463976000|Morning Reports|||0|0||A full round-up of news, sport and business for the day ahead, and a look at the morning's newspapers.(r)
BBC Radio 5 live|1463976900|Wake Up to Money|||0|0||Sean Farrington and Mickey Clark present financial news stories.(r)
BBC Radio 5 live|1463979600|5 Live Breakfast|||0|0||Nicky Campbell and Clare McDonnell present news from the UK and around the world, including business, travel updates and the day's sports stories. Plus, a phone-in on the big issue of the day at 9.00.(r)
BBC Radio 5 live|1463994000|5 Live Daily|||0|0||Adrian Chiles presents news and current affairs interviews. Plus, listeners' stories and contributions, and a round-up of the day's headlines.(r)
BBC Radio 5 live|1464004800|Afternoon Edition|||0|0||Sarah Brett and Adil Ray present an afternoon of engaging stories and conversation, including the latest from the day's news. Featuring big-name interviews, and experts with advice on the latest in health, gadgets, science and media.(r)
BBC Radio 5 live|1464015600|5 Live Drive|||0|0||News, sport and travel updates, with Anna Foster and Tony Livesey.(r)
BBC Radio 5 live|1464026400|5 Live Sport: The Monday Night Club|||0|0||Mark Chapman introduces a football debate following the weekend's cup and international action, with panellists including Robbie Savage and Jonathan Northcroft.
BBC Radio 5 live|1464033600|5 Live Sport: The Tuffers and Vaughan Cricket Show|||0|0||Michael Vaughan and Phil Tufnell discuss cricketing issues, following events at Headingley in the First Test between England and Sri Lanka.
BBC Radio 5 live|1464039000|Phil Williams|||0|0||Dotun Adebayo sits in for Phil Williams with live news and sport. Plus, listeners' emails, texts and tweets.(r)
BBC Radio 5 live|1464048000|Up All Night|||0|0||Rhod Sharp presents stories from around the world. Including an exploration of the frontiers of the web in Outriders and archaeology with Win Scutt.(n)
BBC Radio 5 live|1464062400|Morning Reports|||0|0||A full round-up of news, sport and business for the day ahead, and a look at the morning's newspapers.(n)
BBC Radio 5 live|1464063300|Wake Up to Money|||0|0||Sean Farrington and Louise Cooper present financial news stories.(n)
BBC Radio 5 live|1464066000|5 Live Breakfast|||0|0||Nicky Campbell and Clare McDonnell present news from the UK and around the world, including business, travel updates and the day's sports stories. Plus, a phone-in on the big issue of the day at 9.00.(n)
BBC Radio 5 live|1464080400|5 Live Daily|||0|0||Adrian Chiles presents news and current affairs interviews. Plus, listeners' stories and contributions, and a round-up of the day's headlines.(n)
BBC Radio 5 live|1464091200|Afternoon Edition|||0|0||Sarah Brett and Adil Ray present an afternoon of engaging stories and conversation, including the latest from the day's news. Featuring big-name interviews, and experts with advice on the latest in health, gadgets, science and media.(n)
BBC Radio 5 live|1464102000|5 Live Drive|||0|0||News, sport and travel updates, with Sima Kotecha and Tony Livesey.(n)
BBC Radio 5 live|1464112800|5 Live Sport|||0|0||Will Perry presents the day's sports news, features and interviews.(n)
BBC Radio 5 live|1464114600|5 Live Sport: 5 Live Tennis|||0|0||Russell Fuller presents tennis news and reaction to today's play at the French Open.(n)
BBC Radio 5 live|1464118200|5 Live Sport|||0|0||Eleanor Oldroyd hears first-hand accounts of survivors of abuse in sport - what happened to them, how they lived through it and how they are dealing with the repercussions.(n)
BBC Radio 5 live|1464125400|Phil Williams|||0|0||Dotun Adebayo sits in for Phil Williams with live news and sport. Plus, listeners' emails, texts and tweets.(n)
BBC Radio 5 live sports extra|1463893200|Coming Up on 5 Live Sports Extra|||0|0||Future broadcasts on the station.(c)
BBC Radio 5 live sports extra|1463910900|Cricket|||0|0||Live ball-by-ball commentary from the County Championship as Lancashire face Surrey.(c)
BBC Radio 5 live sports extra|1463929200|Swimming: European Championships|||0|0||Live coverage of the European Swimming Championships as the London Aquatic Centre.(c)
BBC Radio 5 live sports extra|1463938200|Coming Up on 5 Live Sports Extra|||0|0||Future broadcasts on the station.(c)
BBC Radio 5 live sports extra|1463979600|Coming Up on 5 Live Sports Extra|||0|0||Future broadcasts on the station.(c)
BBC Radio 5 live sports extra|1463997300|Cricket|||0|0||Live ball-by-ball commentary from the County Championship as Lancashire face Surrey.(c)
BBC Radio 5 live sports extra|1464024600|Coming Up on 5 Live Sports Extra|||0|0||Future broadcasts on the station.(c)
BBC Radio 5 live sports extra|1464066000|Coming Up on 5 Live Sports Extra|||0|0||Future broadcasts on the station.(n)
BBC Radio 5 live sports extra|1464083700|Cricket|||0|0||Live ball-by-ball commentary from the County Championship as Lancashire face Surrey.(n)
BBC Radio 5 live sports extra|1464111000|Coming Up on 5 Live Sports Extra|||0|0||Future broadcasts on the station.(n)
BBC Radio 6 Music|1463871600|Stuart Maconie's Freakier Zone|||0|0||Musical rarities.(r)
BBC Radio 6 Music|1463875200|The Joy of 6|||0|0||A chance to catch up with the best interviews and moments from the past week on 6 Music.(r)
BBC Radio 6 Music|1463878800|6 Music Recommends|||0|0||The best of the releases featured on Roundtable.(r)
BBC Radio 6 Music|1463882400|6 Music Live Hour|||0|0||Crashland at Cardiff University in 2000, plus archive BBC sessions by Mac DeMarco and Pink Kross. Presented by Chris Hawkins.(r)
BBC Radio 6 Music|1463886000|Race with the Devil: The Gene Vincent Story|||0|0||Roger Daltrey presents profile of rock 'n' roll singer Gene Vincent, who struggled to maintain the early promise of his first hit Be-Bop-a-Lula and moved to England in 1963, where he influenced the style of Lennon and McCartney, Ray Davies, Pete Townshend and Eric Burdon. The programmes features extracts from the play Be-Bop-a-Lula by Rex Weiner about Vincent's friendship with tour mate Eddie Cochrane, who died in a crash in 1960. Part of the Fifties Season.
BBC Radio 6 Music|1463889600|Chris Hawkins|||0|0||Music and chat.(r)
BBC Radio 6 Music|1463896800|Mary Anne Hobbs|||0|0||The DJ presents new music and classic songs.(r)
BBC Radio 6 Music|1463907600|Cerys on 6|||0|0||Eclectic music, poetry and live sessions, presented by former Catatonia singer Cerys Matthews.(r)
BBC Radio 6 Music|1463918400|New Rose and 40 Years of The Damned|||0|0||
BBC Radio 6 Music|1463922000|Guy Garvey's Finest Hour|||0|0||Guests, music and showbiz tales with the Elbow frontman.(r)
BBC Radio 6 Music|1463929200|John Grant's Sunday Service|||0|0||The American singer-songwriter sits in for Jarvis Cocker.(r)
BBC Radio 6 Music|1463936400|Now Playing @6Music|||0|0||Tom Robinson presents a show aiming to provide 6 Music listeners and the online music community with an outlet to recommend, curate and share music.(r)
BBC Radio 6 Music|1463943600|Stuart Maconie's Freak Zone|||0|0||Musical rarities, weird requests and listeners' demos.(r)
BBC Radio 6 Music|1463950800|Don Letts|||0|0||The usual eclectic mix of music and this week's Crucial Vinyl is Aswad's Showcase, which was released in 1981.(r)
BBC Radio 6 Music|1463958000|Guy Garvey's Finest Hour|||0|0||Guests, music and showbiz tales with the Elbow frontman.(r)
BBC Radio 6 Music|1463965200|The BBC Introducing Mixtape|||0|0||Tom Robinson presents a selection of tracks from BBC Introducing.(r)
BBC Radio 6 Music|1463968800|6 Music Live Hour|||0|0||Wildlife at the BBC's Paris Theatre in 1980, plus archive sessions by Zero 7 and Malka Spigel. Presented by Chris Hawkins.(r)
BBC Radio 6 Music|1463972400|Legends of the Dance Floor - A Piece of Paradise|||0|0||Eddie Gordon celebrates the influence of the Paradise Garage nightclub, which operated from 1976 to 1987 in Manhattan and was the base for pioneering DJ Larry Levan. First aired in 2011.(r)
BBC Radio 6 Music|1463976000|Chris Hawkins|||0|0||Music and chat.(r)
BBC Radio 6 Music|1463983200|Nemone|||0|0||Sitting in for Shaun Keaveny.(r)
BBC Radio 6 Music|1463994000|Lauren Laverne|||0|0||New music, live sessions, archive tracks and chat.(r)
BBC Radio 6 Music|1464004800|Mark Radcliffe and Stuart Maconie|||0|0||Tony Parsons chats to Mark and Stuart about his new thriller The Slaughter Man, the latest in his series featuring detective Max Wolfe.(r)
BBC Radio 6 Music|1464015600|Tom Ravenscroft|||0|0||Sitting in for Steve Lamacq.(r)
BBC Radio 6 Music|1464026400|Marc Riley|||0|0||With a live session by Cardiff-based singer-songwriter Cate Le Bon, whose latest album Crab Day was released last month.(r)
BBC Radio 6 Music|1464033600|Gideon Coe|||0|0||The host introduces selected recordings, John Peel sessions and concerts from the BBC archive by a variety of bands past and present.(r)
BBC Radio 6 Music|1464044400|6 Music Recommends|||0|0||The DJ curates an hour of her favourite new releases, showcasing musical genres from folk to hip-hop and African music to electronica.(n)
BBC Radio 6 Music|1464048000|Legends of the Dance Floor - A Piece of Paradise|||0|0||Eddie Gordon continues his documentary celebrating the Paradise Garage nightclub and DJ Larry Levan.(n)
BBC Radio 6 Music|1464051600|Choo Choo Ch'Boogie: The Louis Jordan Story|||0|0||The Wire star Clarke Peters tells the story of the bandleader and musician whose songs bridged the gap between the swing era and R'n'B. Songwriter Jesse Stone is among those recalling the stories behind songs such as Caldonia, Saturday Night Fish Fry, Ain't Nobody Here But Us Chickens. Plus, the inside story of the smash hit Five Guys Named Moe based on Jordan's life, written by and starring Clarke.(n)
BBC Radio 6 Music|1464053400|6 Music Live Hour|||0|0||Robyn Hitchcock & the Egyptians at London's Town & Country Club in 1991, plus archive BBC sessions by Mudhoney and Oasis. Presented by Chris Hawkins.(n)
BBC Radio 6 Music|1464057000|6 Music's Jukebox|||0|0||New tracks, sessions and indie classics.(n)
BBC Radio 6 Music|1464062400|Chris Hawkins|||0|0||Music and chat.(n)
BBC Radio 6 Music|1464069600|Nemone|||0|0||Guests, features and listeners' requests.(n)
BBC Radio 6 Music|1464080400|Lauren Laverne|||0|0||New music, live sessions, archive tracks and chat.(n)
BBC Radio 6 Music|1464091200|Mark Radcliffe and Stuart Maconie|||0|0||Singer-songwriter Graham Nash chats to Shaun about his latest album This Path Tonight, his first solo record for 14 years.(n)
BBC Radio 6 Music|1464102000|Tom Ravenscroft|||0|0||Sitting in for Steve Lamacq.(n)
BBC Radio 6 Music|1464112800|Marc Riley|||0|0||With a live session by Falkirk singer-songwriter Malcolm Middleton, whose new album Summer of '13 is released on Friday.(n)
BBC Radio 6 Music|1464120000|Gideon Coe|||0|0||The host introduces selected recordings, John Peel sessions and concerts from the BBC archive by a variety of bands past and present.(n)
BBC Radio 1Xtra|1463875200|DJ Target|||0|0||The home of new talent.(r)
BBC Radio 1Xtra|1463886000|Diplo and Friends|||0|0||Dance music.(r)
BBC Radio 1Xtra|1463893200|Ace|||0|0||Music, chat and listeners' requests.(r)
BBC Radio 1Xtra|1463907600|Nick Bright|||0|0||Music and chat.(r)
BBC Radio 1Xtra|1463918400|Jamz Supernova|||0|0||The best in new and upfront R'n'B.(r)
BBC Radio 1Xtra|1463929200|DJ Target|||0|0||The home of new talent.(r)
BBC Radio 1Xtra|1463940000|David Rodigan|||0|0||The DJ showcases his love of reggae, playing a selection of classic tunes accompanied by stories from the genre's history.(r)
BBC Radio 1Xtra|1463947200|BBC Radio 1 and 1Xtra's Stories|||0|0||
BBC Radio 1Xtra|1463950800|DJ Edu - Destination Africa|||0|0||The best new underground music from the continent - from hip-hop and R'n'B to afrobeats and azonto.(r)
BBC Radio 1Xtra|1463961600|Monki|||0|0||Music from all corners of the club, featuring house and grime.(r)
BBC Radio 1Xtra|1463972400|DJ Edu - Destination Africa|||0|0||The best new underground music from the continent - from hip-hop and R'n'B to afrobeats and azonto.(r)
BBC Radio 1Xtra|1463983200|Twin B and Yasmin Evans|||0|0||The Breakfast Show.(r)
BBC Radio 1Xtra|1463994000|Trevor Nelson|||0|0||With music from 1Xtra's Live Lounge. Plus, the latest 1Xtra News at 12pm.(r)
BBC Radio 1Xtra|1464003900|Newsbeat|||0|0||Headlines from around the world.(r)
BBC Radio 1Xtra|1464004800|A.Dot|||0|0||Rapper Amplify Dot offers a weekly wrap-up of events and sounds.(r)
BBC Radio 1Xtra|1464015600|Charlie Sloth|||0|0||Hip-hop and heavy hits.(r)
BBC Radio 1Xtra|1464021900|Newsbeat|||0|0||Headlines from around the world.(r)
BBC Radio 1Xtra|1464022800|Charlie Sloth|||0|0||Hip-hop and heavy hits.(r)
BBC Radio 1Xtra|1464026400|MistaJam|||0|0||The DJ plays dubstep, funky, grime, hip-hop, R'n'B, drum 'n' bass, house and dancehall.(r)
BBC Radio 1Xtra|1464037200|Monki|||0|0||Music from all corners of the club, featuring house and grime.(r)
BBC Radio 1Xtra|1464048000|Friction|||0|0||Drum 'n' bass.(n)
BBC Radio 1Xtra|1464058800|Friction|||0|0||Drum 'n' bass.(n)
BBC Radio 1Xtra|1464069600|Twin B and Yasmin Evans|||0|0||The Breakfast Show.(n)
BBC Radio 1Xtra|1464080400|Trevor Nelson|||0|0||With music from 1Xtra's Live Lounge. Plus, the latest 1Xtra News at 12pm.(n)
BBC Radio 1Xtra|1464090300|Newsbeat|||0|0||Headlines from around the world.(n)
BBC Radio 1Xtra|1464091200|A.Dot|||0|0||Rapper Amplify Dot offers a weekly wrap-up of events and sounds.(n)
BBC Radio 1Xtra|1464102000|Charlie Sloth|||0|0||Hip-hop and heavy hits.(n)
BBC Radio 1Xtra|1464108300|Newsbeat|||0|0||Headlines from around the world.(n)
BBC Radio 1Xtra|1464109200|Charlie Sloth|||0|0||Hip-hop and heavy hits.(n)
BBC Radio 1Xtra|1464112800|MistaJam|||0|0||The DJ plays dubstep, funky, grime, hip-hop, R'n'B, drum 'n' bass, house and dancehall.(n)
BBC Radio 1Xtra|1464123600|Jamz Supernova|||0|0||The best in new and upfront R'n'B.(n)
BBC World Service|1463871600|News|||0|0||
BBC World Service|1463871960|The World This Week|||0|0||
BBC World Service|1463873400|The Conversation|||0|0||
BBC World Service|1463875200|News|||0|0||
BBC World Service|1463875560|The Newsroom|||0|0||
BBC World Service|1463876400|Sports News|||0|0||
BBC World Service|1463877000|Outlook|||0|0||Perspectives on important issues.(r)
BBC World Service|1463878800|News|||0|0||
BBC World Service|1463879160|The History Hour|||0|0||
BBC World Service|1463882400|News|||0|0||
BBC World Service|1463882760|Global Business|||0|0||The latest news from the business world.(r)
BBC World Service|1463884200|Heart and Soul|||0|0||The world's main faiths and the personal side of religious belief.(r)
BBC World Service|1463886000|News|||0|0||
BBC World Service|1463886360|The Documentary|||0|0||Investigating global developments, issues and affairs.(r)
BBC World Service|1463889600|News|||0|0||
BBC World Service|1463889960|The Inquiry|||0|0||
BBC World Service|1463891400|The Cultural Frontline|||0|0||
BBC World Service|1463893200|Weekend|||0|0||
BBC World Service|1463902200|Outlook|||0|0||Perspectives on important issues.(r)
BBC World Service|1463904000|News|||0|0||
BBC World Service|1463904360|From Our Own Correspondent|||0|0||Global reports as BBC correspondents across the world tell stories and examine news developments in their region.(r)
BBC World Service|1463905800|Heart and Soul|||0|0||The world's main faiths and the personal side of religious belief.(r)
BBC World Service|1463907600|News|||0|0||
BBC World Service|1463907960|The Compass|||0|0||
BBC World Service|1463909400|Trending|||0|0||
BBC World Service|1463910600|Over to You|||0|0||A chance for listeners to provide feedback on World Service programmes.(r)
BBC World Service|1463911200|News|||0|0||
BBC World Service|1463911560|Global Business|||0|0||The latest news from the business world.(r)
BBC World Service|1463913000|Boston Calling|||0|0||The news from an American perspective.(r)
BBC World Service|1463914800|News|||0|0||
BBC World Service|1463915160|World Questions|||0|0||
BBC World Service|1463918400|Newshour|||0|0||The stories behind the latest headlines.(r)
BBC World Service|1463922000|News|||0|0||
BBC World Service|1463922360|The Documentary|||0|0||Investigating global developments, issues and affairs.(r)
BBC World Service|1463925600|News|||0|0||
BBC World Service|1463925960|The Arts Hour|||0|0||
BBC World Service|1463929200|News|||0|0||
BBC World Service|1463929560|Sportsworld|||0|0||Reports, interviews and analysis.(r)
BBC World Service|1463932800|News|||0|0||
BBC World Service|1463933160|Sportsworld|||0|0||Reports, interviews and analysis.(r)
BBC World Service|1463936400|News|||0|0||
BBC World Service|1463936760|Sportsworld|||0|0||Reports, interviews and analysis.(r)
BBC World Service|1463940000|The Newsroom|||0|0||
BBC World Service|1463941800|Heart and Soul|||0|0||The world's main faiths and the personal side of religious belief.(r)
BBC World Service|1463943600|News|||0|0||
BBC World Service|1463943960|Global Beats|||0|0||
BBC World Service|1463947200|Newshour|||0|0||The stories behind the latest headlines.(r)
BBC World Service|1463950800|News|||0|0||
BBC World Service|1463951160|The History Hour|||0|0||
BBC World Service|1463954400|News|||0|0||
BBC World Service|1463954760|From Our Own Correspondent|||0|0||Global reports as BBC correspondents across the world tell stories and examine news developments in their region.(r)
BBC World Service|1463956200|Global Business|||0|0||The latest news from the business world.(r)
BBC World Service|1463958000|The Newsroom|||0|0||
BBC World Service|1463959200|Sports News|||0|0||The latest stories and results from around the world.(r)
BBC World Service|1463959800|Boston Calling|||0|0||The news from an American perspective.(r)
BBC World Service|1463961600|News|||0|0||
BBC World Service|1463961960|World Business Report|||0|0||Financial news.(r)
BBC World Service|1463963400|The Food Chain|||0|0||
BBC World Service|1463965200|News|||0|0||
BBC World Service|1463965560|The Forum|||0|0||Bridget Kendall invites experts in their respective fields to engage in thought-provoking discussion on a range of topics.(r)
BBC World Service|1463968200|Over to You|||0|0||A chance for listeners to provide feedback on World Service programmes.(r)
BBC World Service|1463968800|News|||0|0||
BBC World Service|1463969160|HARDtalk|||0|0||Interviews with newsmakers and personalities from across the globe.(r)
BBC World Service|1463970600|The Why Factor|||0|0||The extraordinary and hidden histories behind everyday objects and actions.(r)
BBC World Service|1463971800|More or Less|||0|0||
BBC World Service|1463972400|News|||0|0||
BBC World Service|1463972760|Newsday|||0|0||The latest headlines.(r)
BBC World Service|1463976000|Newsday|||0|0||The latest headlines.(r)
BBC World Service|1463977800|The Conversation|||0|0||
BBC World Service|1463979600|Newsday|||0|0||The latest headlines.(r)
BBC World Service|1463988600|Business Daily|||0|0||Business and finance news, interviews and reports.(r)
BBC World Service|1463989800|Witness|||0|0||
BBC World Service|1463990400|News|||0|0||
BBC World Service|1463990760|The Arts Hour|||0|0||
BBC World Service|1463994000|World Update|||0|0||
BBC World Service|1463997600|Outside Source|||0|0||
BBC World Service|1464001200|News|||0|0||
BBC World Service|1464001560|Outlook|||0|0||Perspectives on important issues.(r)
BBC World Service|1464004800|The Newsroom|||0|0||
BBC World Service|1464006600|The Conversation|||0|0||
BBC World Service|1464008400|Newshour|||0|0||The stories behind the latest headlines.(r)
BBC World Service|1464012000|News|||0|0||
BBC World Service|1464012360|HARDtalk|||0|0||Interviews with newsmakers and personalities from across the globe.(r)
BBC World Service|1464013800|The Why Factor|||0|0||The extraordinary and hidden histories behind everyday objects and actions.(r)
BBC World Service|1464015000|More or Less|||0|0||
BBC World Service|1464015600|News|||0|0||
BBC World Service|1464015960|Business Daily|||0|0||Business and finance news, interviews and reports.(r)
BBC World Service|1464017100|The Essential: Trending|||0|0||
BBC World Service|1464017400|Sport Today|||0|0||News and results from around the world.(r)
BBC World Service|1464019200|World Have Your Say|||0|0||
BBC World Service|1464022800|The Newsroom|||0|0||
BBC World Service|1464024600|World Business Report|||0|0||Financial news.(r)
BBC World Service|1464026400|The Newsroom|||0|0||
BBC World Service|1464028200|The Conversation|||0|0||
BBC World Service|1464030000|News|||0|0||
BBC World Service|1464030360|Outlook|||0|0||Perspectives on important issues.(r)
BBC World Service|1464033600|Newshour|||0|0||The stories behind the latest headlines.(r)
BBC World Service|1464037200|News|||0|0||
BBC World Service|1464037560|HARDtalk|||0|0||Interviews with newsmakers and personalities from across the globe.(r)
BBC World Service|1464039000|Discovery|||0|0||Insights from leading scientific figures.(r)
BBC World Service|1464040800|The Newsroom|||0|0||
BBC World Service|1464042000|Sports News|||0|0||
BBC World Service|1464042600|World Business Report|||0|0||Financial news.(r)
BBC World Service|1464044400|News|||0|0||
BBC World Service|1464044760|The Arts Hour|||0|0||
BBC World Service|1464048000|News|||0|0||
BBC World Service|1464048360|Business Matters|||0|0||
BBC World Service|1464051600|News|||0|0||
BBC World Service|1464051960|Outlook|||0|0||Perspectives on important issues.(n)
BBC World Service|1464055200|News|||0|0||
BBC World Service|1464055560|The Inquiry|||0|0||
BBC World Service|1464057000|Discovery|||0|0||Insights from leading scientific figures.(n)
BBC World Service|1464058800|Newsday|||0|0||The latest headlines.(n)
BBC World Service|1464062400|Newsday|||0|0||The latest headlines.(n)
BBC World Service|1464064200|The Documentary|||0|0||Investigating global developments, issues and affairs.(n)
BBC World Service|1464066000|Newsday|||0|0||The latest headlines.(n)
BBC World Service|1464075000|Business Daily|||0|0||Business and finance news, interviews and reports.(n)
BBC World Service|1464076200|Witness|||0|0||
BBC World Service|1464076800|News|||0|0||
BBC World Service|1464077160|The Forum|||0|0||Bridget Kendall invites experts in their respective fields to engage in thought-provoking discussion on a range of topics.(n)
BBC World Service|1464079800|Sporting Witness|||0|0||
BBC World Service|1464080400|World Update|||0|0||
BBC World Service|1464084000|Outside Source|||0|0||
BBC World Service|1464087600|News|||0|0||
BBC World Service|1464087960|Outlook|||0|0||Perspectives on important issues.(n)
BBC World Service|1464091200|The Newsroom|||0|0||
BBC World Service|1464093000|The Documentary|||0|0||Investigating global developments, issues and affairs.(n)
BBC World Service|1464094800|Newshour|||0|0||The stories behind the latest headlines.(n)
BBC World Service|1464098400|News|||0|0||
BBC World Service|1464098760|The Inquiry|||0|0||
BBC World Service|1464100200|Discovery|||0|0||Insights from leading scientific figures.(n)
BBC World Service|1464102000|News|||0|0||
BBC World Service|1464102360|Business Daily|||0|0||Business and finance news, interviews and reports.(n)
BBC World Service|1464103500|The Essential|||0|0||
BBC World Service|1464103800|Sport Today|||0|0||News and results from around the world.(n)
BBC World Service|1464105600|World Have Your Say|||0|0||
BBC World Service|1464109200|The Newsroom|||0|0||
BBC World Service|1464111000|World Business Report|||0|0||Financial news.(n)
BBC World Service|1464112800|The Newsroom|||0|0||
BBC World Service|1464114600|The Documentary|||0|0||Investigating global developments, issues and affairs.(n)
BBC World Service|1464116400|News|||0|0||
BBC World Service|1464116760|Outlook|||0|0||Perspectives on important issues.(n)
BBC World Service|1464120000|Newshour|||0|0||The stories behind the latest headlines.(n)
BBC World Service|1464123600|News|||0|0||
BBC World Service|1464123960|The Inquiry|||0|0||
BBC World Service|1464125400|Click|||0|0||Technological and digital news from around the world.(n)
BBC World Service|1464127200|The Newsroom|||0|0||
BBC World Service|1464128400|Sports News|||0|0||
BBC World Service|1464129000|World Business Report|||0|0||Financial news.(n)
BBC Asian Network|1463871600|As Radio 5 Live|||0|0||
BBC Asian Network|1463893200|Harpz Kaur|||0|0||
BBC Asian Network|1463907600|Gagan Grewal|||0|0||News, music and features.(r)
BBC Asian Network|1463918400|Asian Network Presents|||0|0||
BBC Asian Network|1463922000|Ashanti Omkar|||0|0||
BBC Asian Network|1463929200|Saima Ajram|||0|0||With Pakistani music and features.(r)
BBC Asian Network|1463936400|Dipps Bhamrah|||0|0||With Bhangra music and Punjabi-based features.(r)
BBC Asian Network|1463943600|Nadia Ali|||0|0||With Bengali music and features.(r)
BBC Asian Network|1463950800|Alpa Pandya|||0|0||Alpa brings the best in Bollywood and Gujarati music, culture and news.(r)
BBC Asian Network|1463958000|As Radio 5 Live|||0|0||
BBC Asian Network|1463979600|Tommy Sandhu|||0|0||The DJ presents lively chat, celebrity guests, the latest headlines and sporting news, along with Bollywood and Bhangra hits.(r)
BBC Asian Network|1463994000|Nihal|||0|0||Topical discussion and debate.(r)
BBC Asian Network|1464004800|Asian Network Reports|||0|0||Hard-hitting documentary.(r)
BBC Asian Network|1464006600|Noreen Khan|||0|0||Lively mix of news, music and chat.(r)
BBC Asian Network|1464019200|Asian Network Reports|||0|0||Hard-hitting documentary.(r)
BBC Asian Network|1464021000|Bobby Friction|||0|0||Cutting-edge British Asian music.(r)
BBC Asian Network|1464033600|Ray Khan|||0|0||
BBC Asian Network|1464044400|As Radio 5 Live|||0|0||
BBC Asian Network|1464066000|Tommy Sandhu|||0|0||The DJ presents lively chat, celebrity guests, the latest headlines and sporting news, along with Bollywood and Bhangra hits.(n)
BBC Asian Network|1464080400|Nihal|||0|0||Topical discussion and debate.(n)
BBC Asian Network|1464091200|Asian Network Reports|||0|0||Hard-hitting documentary.(n)
BBC Asian Network|1464093000|Noreen Khan|||0|0||Lively mix of news, music and chat.(n)
BBC Asian Network|1464105600|Asian Network Reports|||0|0||Hard-hitting documentary.(n)
BBC Asian Network|1464107400|Bobby Friction|||0|0||Cutting-edge British Asian music.(n)
BBC Asian Network|1464120000|Ray Khan|||0|0||
