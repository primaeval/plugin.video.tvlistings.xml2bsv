BBC One|BBC1|http://my.tvguide.co.uk/channel_logos/70.png|000000=
BBC Two|BBC2|http://my.tvguide.co.uk/channel_logos/89.png|000001=
BBC Four|BBC4|http://my.tvguide.co.uk/channel_logos/109.png|000002=
CBBC|CBBC|http://my.tvguide.co.uk/channel_logos/118.png|000003=
CBeebies|CBeebies|http://my.tvguide.co.uk/channel_logos/119.png|000004=
BBC News|BBC News|http://my.tvguide.co.uk/channel_logos/66.png|000005=
BBC Parliament|BBC Parliament|http://my.tvguide.co.uk/channel_logos/67.png|000006=
Channel 4|Channel 4|http://my.tvguide.co.uk/channel_logos/121.png|000007=
More4|More4|http://my.tvguide.co.uk/channel_logos/361.png|000008=
Film4|Film4|http://my.tvguide.co.uk/channel_logos/145.png|000009=
ITV Anglia|ITV Anglia|http://my.tvguide.co.uk/channel_logos/165.png|000010=
ITV2|ITV2|http://my.tvguide.co.uk/channel_logos/180.png|000011=
ITV3|ITV3|http://my.tvguide.co.uk/channel_logos/360.png|000012=
ITV4|ITV4|http://my.tvguide.co.uk/channel_logos/367.png|000013=
CITV|CITV|http://my.tvguide.co.uk/channel_logos/382.png|000014=
Channel 5|Channel 5|http://my.tvguide.co.uk/channel_logos/148.png|000015=
Sky Sports 1|Sky Sports 1|http://my.tvguide.co.uk/channel_logos/260.png|000016=
Sky Sports 2|Sky Sports 2|http://my.tvguide.co.uk/channel_logos/261.png|000017=
Sky Sports 3|Sky Sports 3|http://my.tvguide.co.uk/channel_logos/262.png|000018=
Sky Sports 4|Sky Sports 4|http://my.tvguide.co.uk/channel_logos/264.png|000019=
Sky Sports 5|Sky Sports 5|http://my.tvguide.co.uk/channel_logos/918.png|000020=
Sky Sports F1|Sky Sports F1|http://my.tvguide.co.uk/channel_logos/736.png|000021=
DR1|DR1||000022=
DR Ramasjang|DRRAMA||000023=
BBC Red Button 1|BBC Red Button 1|http://my.tvguide.co.uk/channel_logos/636.png|000024=
BBC Red Button 2|BBC Red Button 2|http://my.tvguide.co.uk/channel_logos/840.png|000025=
BBC Red Button 3|BBC Red Button 3|http://my.tvguide.co.uk/channel_logos/767.png|000026=
BBC Red Button 4|BBC Red Button 4|http://my.tvguide.co.uk/channel_logos/914.png|000027=
BBC Red Button 5|BBC Red Button 5|http://my.tvguide.co.uk/channel_logos/915.png|000028=
BBC Red Button HD|BBC Red Button HD|http://my.tvguide.co.uk/channel_logos/766.png|000029=
BBC Sport Interactive BBC1|BBC Sport Interactive BBC1|http://my.tvguide.co.uk/channel_logos/643.png|000030=
BBC Sport Interactive BBC2|BBC Sport Interactive BBC2|http://my.tvguide.co.uk/channel_logos/644.png|000031=
BBC Sport Interactive BBC3|BBC Sport Interactive BBC3|http://my.tvguide.co.uk/channel_logos/651.png|000032=
BBC Radio 1|BBC Radio 1||000033=
BBC Radio 2|BBC Radio 2||000034=
BBC Radio 3|BBC Radio 3||000035=
BBC Radio 4 FM|BBC Radio 4 FM||000036=
BBC Radio 4 Extra|BBC Radio 4 Extra||000037=
BBC Radio 4 LW|BBC Radio 4 LW||000038=
BBC Radio 5 live|BBC Radio 5 live||000039=
BBC Radio 5 live sports extra|BBC Radio 5 live sports extra||000040=
BBC Radio 6 Music|BBC Radio 6 Music||000041=
BBC Radio 1Xtra|BBC Radio 1Xtra||000042=
BBC World Service|BBC World Service||000043=
BBC Asian Network|BBC Asian Network||000044=
